* AND Gate
.include /data/yaohuihan/Research/STA_Modeling/Spice/Libs/FreePDK/subckts/AND2X1.pex.netlist
.include /data/yaohuihan/Research/STA_Modeling/Spice/Libs/FreePDK/subckts/AND2X1.pex.netlist.AND2X1.pxi
.include /data/yaohuihan/Research/STA_Modeling/Spice/Libs/FreePDK/gpdk45nm.m

.temp 27
.param VOL=1.1
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 1.35000n 1.35000n 50n 500n)
VIN_B b 0 DC VOL

Cout y 0 0.20000p

X1 y an b VDD VSS AND2X1

.tran 0.000001n 300n

.measure tran tpHL TRIG V(an) VAL=0.55 FALL=1 TARG V(y) VAL=0.55 FALL=1
.measure tran tpLH TRIG V(an) VAL=0.55 RISE=1 TARG V(y) VAL=0.55 RISE=1

.end
