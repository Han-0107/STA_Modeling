* NAND Gate
.include ./Libs/cells.sp
.include ./Libs/gpdk45nm.m

.param VOL=3
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 2.0n 2.0n 20n 40n)
VIN_B b 0 DC VOL

Cout y 0 0.2p

X1 y an b VDD VSS NAND2X1

.tran 0.0001n 25n

.control
run
meas tran tpHL TRIG V(an) VAL=2.5 FALL=1 TARG V(y) VAL=2.5 RISE=1
meas tran tpLH TRIG V(an) VAL=2.5 RISE=1 TARG V(y) VAL=2.5 FALL=1

echo "tpHL = " $&tpHL > ./Delays/nand_VOL_nand_VOL_3_Trans_2.0n_Cap_0.2p.txt.txt
echo "tpLH = " $&tpLH >> ./Delays/nand_VOL_nand_VOL_3_Trans_2.0n_Cap_0.2p.txt.txt
.endc

.end
