* NOT Gate
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/FreePDK/cells.sp
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/FreePDK/gpdk45nm.m

.temp 27
.param VOL=1.1
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 0.1n 0.1n 5n 40n)

Cout y 0 0.1p

X1 y an VDD VSS INVX1

.tran 0.000001n 10n

.measure tran tpHL TRIG V(an) VAL=0.55 FALL=1 TARG V(y) VAL=0.55 RISE=1
.measure tran tpLH TRIG V(an) VAL=0.55 RISE=1 TARG V(y) VAL=0.55 FALL=1

.end
