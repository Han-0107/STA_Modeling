* NAND Gate
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/FreePDK/cells.sp
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/FreePDK/gpdk45nm.m

.temp 27
.param VOL=1.2
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 0.40000n 0.40000n 50n 500n)
VIN_B b 0 DC VOL

Cout y 0 5.00000p

X1 y an b VDD VSS NAND2X1

.tran 0.000001n 300n

.measure tran tpHL TRIG V(an) VAL=0.6 FALL=1 TARG V(y) VAL=0.6 RISE=1
.measure tran tpLH TRIG V(an) VAL=0.6 RISE=1 TARG V(y) VAL=0.6 FALL=1

.end