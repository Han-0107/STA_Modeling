* AND Gate
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/FreePDK/cells.sp
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/FreePDK/gpdk45nm.m

.temp 27
.param VOL=1.11
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 0.10000n 0.10000n 50n 500n)
VIN_B b 0 DC VOL

Cout y 0 0.10000p

X1 y an b VDD VSS AND2X1

.tran 0.000001n 300n

.measure tran tpHL TRIG V(an) VAL=0.555 FALL=1 TARG V(y) VAL=0.555 FALL=1
.measure tran tpLH TRIG V(an) VAL=0.555 RISE=1 TARG V(y) VAL=0.555 RISE=1

.end
