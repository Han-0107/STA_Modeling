* NAND Gate
.include ./Libs/cells.sp
.include ./Libs/gpdk45nm.m

.param VOL=1.1
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 1n 1n 20n 40n)
VIN_B b 0 DC VOL

Cout y 0 0.1p

X1 y an b VDD VSS NAND2X1

.tran 0.0001n 25n

.control
run
meas tran tpHL TRIG V(an) VAL=0.55 FALL=1 TARG V(y) VAL=0.55 RISE=1
meas tran tpLH TRIG V(an) VAL=0.55 RISE=1 TARG V(y) VAL=0.55 FALL=1

echo "tpHL = " $&tpHL > ./Delays/nand_VOL_1.1V.txt
echo "tpLH = " $&tpLH >> ./Delays/nand_VOL_1.1V.txt
.endc

.end
