***********************************************************************
****                                                               ****
****  The data contained in the file is created for educational    **** 
****  and training purposes only and are not recommended           ****
****  for fabrication                                              ****
****                                                               ****
***********************************************************************
****                                                               ****
****  Copyright (C) 2013 Synopsys, Inc.                            ****
****                                                               ****
***********************************************************************
****                                                               ****
****  The 32/28nm Generic Library ("Library") is unsupported       ****    
****  Confidential Information of Synopsys, Inc. ("Synopsys")      ****    
****  provided to you as Documentation under the terms of the      ****    
****  End User Software License Agreement between you or your      ****    
****  employer and Synopsys ("License Agreement") and you agree    ****    
****  not to distribute or disclose the Library without the        ****    
****  prior written consent of Synopsys. The Library IS NOT an     ****    
****  item of Licensed Software or Licensed Product under the      ****    
****  License Agreement.  Synopsys and/or its licensors own        ****    
****  and shall retain all right, title and interest in and        ****    
****  to the Library and all modifications thereto, including      ****    
****  all intellectual property rights embodied therein. All       ****    
****  rights in and to any Library modifications you make are      ****    
****  hereby assigned to Synopsys. If you do not agree with        ****    
****  this notice, including the disclaimer below, then you        ****    
****  are not authorized to use the Library.                       ****    
****                                                               ****  
****                                                               ****      
****  THIS LIBRARY IS BEING DISTRIBUTED BY SYNOPSYS SOLELY ON AN   ****
****  "AS IS" BASIS, WITH NO INTELLECUTAL PROPERTY                 ****
****  INDEMNIFICATION AND NO SUPPORT. ANY EXPRESS OR IMPLIED       ****
****  WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED       ****
****  WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR   ****
****  PURPOSE ARE HEREBY DISCLAIMED. IN NO EVENT SHALL SYNOPSYS    ****
****  BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     ****
****  EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT      ****
****  LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;     ****
****  LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)     ****
****  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN    ****
****  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE    ****
****  OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS      ****
****  DOCUMENTATION, EVEN IF ADVISED OF THE POSSIBILITY OF         ****
****  SUCH DAMAGE.                                                 **** 		
****                                                               ****  
***********************************************************************




.subckt AND2X1_RVT A1 A2 VDD VSS Y
MN3 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP3 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
.ends AND2X1_RVT




.subckt AND2X2_RVT A1 A2 VDD VSS Y
MP1 Y1 A1 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP3 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP2 Y1 A2 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
.ends AND2X2_RVT




.subckt AND2X4_RVT A1 A2 VDD VSS Y
MP1 Y1 A1 VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MP3 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MN3 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN2 SA1 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends AND2X4_RVT




.subckt AND3X1_RVT A1 A2 A3 VDD VSS Y
MN3 SA2 A3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP3 Y1 A3 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP4 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
.ends AND3X1_RVT




.subckt AND3X2_RVT A1 A2 A3 VDD VSS Y
MP3 Y1 A3 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP4 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP1 Y1 A1 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA2 A3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
.ends AND3X2_RVT




.subckt AND3X4_RVT A1 A2 A3 VDD VSS Y
MP3 Y1 A3 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP4 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MP1 Y1 A1 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA2 A3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
.ends AND3X4_RVT




.subckt AND4X1_RVT A1 A2 A3 A4 VDD VSS Y
MN4 SA3 A4 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN3 SA2 A3 SA3 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP4 Y1 A4 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP5 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP3 Y1 A3 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
.ends AND4X1_RVT




.subckt AND4X2_RVT A1 A2 A3 A4 VDD VSS Y
MP7 Y Y3 VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP6 Y3 Y2 VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP4 Y1 A1 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP3 Y1 A2 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP2 Y1 A3 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP1 Y1 A4 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP5 Y2 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MN7 Y Y3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN6 Y3 Y2 VSS VSS n105 w=0.27u l=0.03u nf=1 m=1
MN2 SA2 A3 SA1 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN3 SA3 A2 SA2 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN5 Y2 Y1 VSS VSS n105 w=0.22u l=0.03u nf=1 m=1
MN4 Y1 A1 SA3 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN1 SA1 A4 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
.ends AND4X2_RVT




.subckt AND4X4_RVT A1 A2 A3 A4 VDD VSS Y
MN7 Y Y3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN6 Y3 Y2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN5 Y2 Y1 VSS VSS n105 w=0.22u l=0.03u nf=1 m=1
MN3 SA3 A2 SA2 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN1 SA1 A4 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN2 SA2 A3 SA1 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN4 Y1 A1 SA3 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MP7 Y Y3 VDD VDD p105 w=0.80u l=0.03u nf=1 m=4
MP6 Y3 Y2 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP5 Y2 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP2 Y1 A3 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP1 Y1 A4 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP4 Y1 A1 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP3 Y1 A2 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
.ends AND4X4_RVT




.subckt ANTENNA_RVT INP VDD VSS
DD7 INP VDD nd area=4p l=2u w=2u m=1
DD6 VSS INP nd area=4p l=2u w=2u m=1
.ends ANTENNA_RVT




.subckt AO21X1_RVT A1 A2 A3 VDD VSS Y
MN2 net3 A1 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN3 net3 A3 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN4 Y net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net2 A2 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MP4 Y net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP2 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP3 net3 A3 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
.ends AO21X1_RVT




.subckt AO21X2_RVT A1 A2 A3 VDD VSS Y
MP1 net1 A2 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP3 net3 A3 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP4 Y net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN1 net2 A2 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN4 Y net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 net3 A3 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN2 net3 A1 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
.ends AO21X2_RVT




.subckt AO221X1_RVT A1 A2 A3 A4 A5 VDD VSS Y
MN2 net5 A1 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN5 net5 A5 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MN6 Y net5 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 net5 A3 net4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net5 A5 net3 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP6 Y net5 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
.ends AO221X1_RVT




.subckt AO221X2_RVT A1 A2 A3 A4 A5 VDD VSS Y
MP1 net1 A2 VDD VDD p105 w=0.67u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.67u l=0.03u nf=1.0 m=1
MP6 Y net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP4 net3 A3 net1 VDD p105 w=0.67u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.67u l=0.03u nf=1.0 m=1
MP5 net5 A5 net3 VDD p105 w=0.67u l=0.03u nf=1.0 m=1
MN4 net5 A3 net4 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN6 Y net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 net5 A5 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN2 net5 A1 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
.ends AO221X2_RVT




.subckt AO222X1_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MP5 net5 A6 net3 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP6 net5 A5 net3 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP7 Y net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MN1 net2 A2 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 net5 A1 net2 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN6 net5 A5 net6 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN4 net5 A3 net4 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN5 net6 A6 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN7 Y net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
.ends AO222X1_RVT




.subckt AO222X2_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MP3 net3 A4 net1 VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP7 Y net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net1 A2 VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 net5 A5 net3 VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP5 net5 A6 net3 VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MN7 Y net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 net6 A6 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN4 net5 A3 net4 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN6 net5 A5 net6 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN2 net5 A1 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
.ends AO222X2_RVT




.subckt AO22X1_RVT A1 A2 A3 A4 VDD VSS Y
MP4 net3 A3 net1 VDD p105 w=0.51u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.51u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.51u l=0.03u nf=1.0 m=1
MP5 Y net3 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.51u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN5 Y net3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net3 A3 net4 VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN2 net3 A1 net2 VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends AO22X1_RVT




.subckt AO22X2_RVT A1 A2 A3 A4 VDD VSS Y
MN1 net2 A2 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN5 Y net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN4 net3 A3 net4 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN2 net3 A1 net2 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.54u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.54u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.54u l=0.03u nf=1.0 m=1
MP5 Y net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP3 net3 A4 net1 VDD p105 w=0.54u l=0.03u nf=1.0 m=1
.ends AO22X2_RVT




.subckt AOBUFX1_RVT A VDD VDDG VSS Y
MN1 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN0 SA1 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP1 Y SA1 VDDG VDDG p105 w=0.8u l=0.03u nf=1.0 m=1
MP0 SA1 A VDDG VDDG p105 w=0.60u l=0.03u nf=1.0 m=1
.ends AOBUFX1_RVT




.subckt AOBUFX2_RVT A VDD VDDG VSS Y
MN1 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN0 SA1 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP1 Y SA1 VDDG VDDG p105 w=0.8u l=0.03u nf=1 m=2
MP0 SA1 A VDDG VDDG p105 w=0.60u l=0.03u nf=1.0 m=1
.ends AOBUFX2_RVT




.subckt AOBUFX4_RVT A VDD VDDG VSS Y
MN1 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN0 SA1 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP1 Y SA1 VDDG VDDG p105 w=0.8u l=0.03u nf=1 m=4
MP0 SA1 A VDDG VDDG p105 w=0.60u l=0.03u nf=1.0 m=1
.ends AOBUFX4_RVT




.subckt AODFFARX1_RVT CLK D Q QN RSTB VDD VDDG VSS
MM19 VDDG net7 net211 VDDG p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net211 net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKN VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDDG VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP26 VDDG net213 net2 VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP14 QN net213 VDDG VDDG p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net2 VDDG VDDG p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net191 D VDDG VDDG p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net7 CLKP net191 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKP VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net213 net2 net4 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP7 net213 CLKN net211 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 net211 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net211 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN25 net3 net213 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN23 net213 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net213 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net191 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net7 CLKN net191 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net213 CLKP net211 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends AODFFARX1_RVT




.subckt AODFFARX2_RVT CLK D Q QN RSTB VDD VDDG VSS
MM19 VDDG net7 net211 VDDG p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net211 net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKN VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDDG VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP26 VDDG net213 net2 VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP14 QN net213 VDDG VDDG p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net2 VDDG VDDG p105 w=0.8u l=0.03u nf=1 m=2
MP01 net191 D VDDG VDDG p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net7 CLKP net191 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKP VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net213 net2 net4 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP7 net213 CLKN net211 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 net211 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net211 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN25 net3 net213 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN23 net213 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net213 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net191 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net7 CLKN net191 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net213 CLKP net211 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends AODFFARX2_RVT




.subckt AODFFNARX1_RVT CLK D Q QN RSTB VDD VDDG VSS
MM19 VDDG net7 net211 VDDG p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net211 net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKP VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDDG VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP26 VDDG net213 net2 VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP14 QN net213 VDDG VDDG p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net2 VDDG VDDG p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net191 D VDDG VDDG p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net7 CLKN net191 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKN VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net213 net2 net4 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP7 net213 CLKP net211 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 net211 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net211 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN25 net3 net213 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN23 net213 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net213 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net191 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net7 CLKP net191 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net213 CLKN net211 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends AODFFNARX1_RVT




.subckt AODFFNARX2_RVT CLK D Q QN RSTB VDD VDDG VSS
MM19 VDDG net7 net211 VDDG p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net211 net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKP VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDDG VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP26 VDDG net213 net2 VDDG p105 w=0.52u l=0.03u nf=1.0 m=1
MP14 QN net213 VDDG VDDG p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net2 VDDG VDDG p105 w=0.8u l=0.03u nf=1 m=2
MP01 net191 D VDDG VDDG p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net7 CLKN net191 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDDG VDDG p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKN VDDG VDDG p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net213 net2 net4 VDDG p105 w=0.3u l=0.03u nf=1 m=1
MP7 net213 CLKP net211 VDDG p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 net211 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net211 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN25 net3 net213 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN23 net213 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net213 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net191 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net7 CLKP net191 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net213 CLKN net211 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends AODFFNARX2_RVT




.subckt AOI21X1_RVT A1 A2 A3 VDD VSS Y
MN5 Y net4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN2 net3 A1 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN3 net3 A3 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN4 net4 net3 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MP5 Y net4 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP4 net4 net3 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP3 net3 A3 net1 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
.ends AOI21X1_RVT




.subckt AOI21X2_RVT A1 A2 A3 VDD VSS Y
MP2 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP3 net3 A3 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP4 net4 net3 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP5 Y net4 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN4 net4 net3 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN3 net3 A3 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN2 net3 A1 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN5 Y net4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
.ends AOI21X2_RVT




.subckt AOI221X1_RVT A1 A2 A3 A4 A5 VDD VSS Y
MN6 net7 net5 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net5 A1 net2 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN5 net5 A5 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN7 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN4 net5 A3 net4 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MP6 net7 net5 VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP5 net5 A5 net3 VDD p105 w=0.54u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP7 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
.ends AOI221X1_RVT




.subckt AOI221X2_RVT A1 A2 A3 A4 A5 VDD VSS Y
MP7 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP3 net3 A4 net1 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP5 net5 A5 net3 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP6 net7 net5 VDD VDD p105 w=0.54u l=0.03u nf=1.0 m=1
MN5 net5 A5 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN4 net5 A3 net4 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN2 net5 A1 net2 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN7 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN6 net7 net5 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
.ends AOI221X2_RVT




.subckt AOI222X1_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MP7 net5 net7 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP8 Y net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP1 net1 A2 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP6 net7 A5 net3 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP5 net7 A6 net3 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MN7 net5 net7 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN8 Y net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN5 net6 A6 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN4 net7 A3 net4 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN3 net4 A4 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN6 net7 A5 net6 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 net7 A1 net2 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
.ends AOI222X1_RVT




.subckt AOI222X2_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MN1 net2 A2 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN4 net7 A3 net4 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN5 net6 A6 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 net7 A1 net2 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN6 net7 A5 net6 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN8 Y net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 net4 A4 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN7 net5 net7 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MP5 net7 A6 net3 VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP8 Y net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP3 net3 A4 net1 VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP6 net7 A5 net3 VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP7 net5 net7 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
.ends AOI222X2_RVT




.subckt AOI22X1_RVT A1 A2 A3 A4 VDD VSS Y
MN5 net4 net3 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 net6 A4 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN6 Y net4 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net3 A3 net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net3 A1 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net4 net3 VDD VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP4 net3 A3 net1 VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP1 net1 A2 VDD VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP6 Y net4 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.53u l=0.03u nf=1.0 m=1
.ends AOI22X1_RVT




.subckt AOI22X2_RVT A1 A2 A3 A4 VDD VSS Y
MP1 net1 A2 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP3 net3 A4 net1 VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP6 Y net4 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP4 net3 A3 net1 VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP2 net1 A1 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP5 net4 net3 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MN4 net3 A3 net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net3 A1 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN6 Y net4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 net6 A4 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net2 A2 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN5 net4 net3 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
.ends AOI22X2_RVT




.subckt AOINVX1_RVT A VDD VDDG VSS Y
MN0 Y A VSS VSS n105 w=0.31u l=0.03u nf=1.0 m=1
MP0 Y A VDDG VDDG p105 w=0.80u l=0.03u nf=1.0 m=1
.ends AOINVX1_RVT




.subckt AOINVX2_RVT A VDD VDDG VSS Y
MN0 Y A VSS VSS n105 w=0.31u l=0.03u nf=1 m=2
MP0 Y A VDDG VDDG p105 w=0.80u l=0.03u nf=1 m=2
.ends AOINVX2_RVT




.subckt AOINVX4_RVT A VDD VDDG VSS Y
MN0 Y A VSS VSS n105 w=0.31u l=0.03u nf=1 m=4
MP0 Y A VDDG VDDG p105 w=0.80u l=0.03u nf=1 m=4
.ends AOINVX4_RVT




.subckt BSLEX1_RVT EN INOUT1 INOUT2 VDD VSS
MN2 INOUT1 EN INOUT2 VSS n105 w=0.375u l=0.03u nf=1.0 m=1
MN1 net35 EN VSS VSS n105 w=0.125u l=0.03u nf=1.0 m=1
MP2 INOUT1 net35 INOUT2 VDD p105 w=0.715u l=0.03u nf=1.0 m=1
MP1 net35 EN VDD VDD p105 w=0.235u l=0.03u nf=1.0 m=1
.ends BSLEX1_RVT




.subckt BSLEX2_RVT EN INOUT1 INOUT2 VDD VSS
MN2 INOUT1 EN INOUT2 VSS n105 w=0.375u l=0.03u nf=1 m=2
MN1 net35 EN VSS VSS n105 w=0.185u l=0.03u nf=1.0 m=1
MP2 INOUT1 net35 INOUT2 VDD p105 w=0.715u l=0.03u nf=1 m=2
MP1 net35 EN VDD VDD p105 w=0.355u l=0.03u nf=1.0 m=1
.ends BSLEX2_RVT




.subckt BSLEX4_RVT EN INOUT1 INOUT2 VDD VSS
MN2 INOUT1 EN INOUT2 VSS n105 w=0.375u l=0.03u nf=1 m=4
MN1 net35 EN VSS VSS n105 w=0.375u l=0.03u nf=1.0 m=1
MP2 INOUT1 net35 INOUT2 VDD p105 w=0.715u l=0.03u nf=1 m=4
MP1 net35 EN VDD VDD p105 w=0.715u l=0.03u nf=1.0 m=1
.ends BSLEX4_RVT




.subckt BUSKP_RVT A VDD VSS
MN5 net194 SA1 net195 VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN4 net192 SA1 net194 VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN3 net190 SA1 net192 VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN2 net188 SA1 net190 VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN1 A SA1 net188 VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN6 net195 SA1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN0 SA1 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP2 A SA1 net185 VDD p105 w=0.20u l=0.03u nf=1.0 m=1
MP1 net185 SA1 VDD VDD p105 w=0.20u l=0.03u nf=1.0 m=1
MP0 SA1 A VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends BUSKP_RVT




.subckt CGLNPRX2_RVT CLK EN GCLK SE VDD VSS
MN7 net75 ENL VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net68 net75 VSS VSS n105 w=0.18u l=0.03u nf=1.0 m=1
MN10 GCLK net68 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN8 net68 CLKP VSS VSS n105 w=0.18u l=0.03u nf=1.0 m=1
MN1 net2 SE VSS VSS n105 w=0.18u l=0.03u nf=1.0 m=1
MN2 net2 EN VSS VSS n105 w=0.18u l=0.03u nf=1.0 m=1
MN11 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN12 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN6 net5 ENL VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 net3 CLKN net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 ENL net3 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 CLKP net3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net75 ENL VDD VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP9 net68 net75 net66 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP10 GCLK net68 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP8 net66 CLKP VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP2 net2 EN net1 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP1 net1 SE VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP5 net4 ENL VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net3 CLKP net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP4 ENL net3 VDD VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP11 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP3 net2 CLKN net3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
.ends CGLNPRX2_RVT




.subckt CGLNPRX8_RVT CLK EN GCLK SE VDD VSS
MP1 net1 SE VDD VDD p105 w=0.75u l=0.03u nf=1.0 m=1
MP3 net2 CLKN net3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net2 EN net1 VDD p105 w=0.75u l=0.03u nf=1.0 m=1
MP12 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP11 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP4 ENL net3 VDD VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP6 net3 CLKP net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP5 net4 ENL VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP8 net13 CLKP VDD VDD p105 w=0.75u l=0.03u nf=1.0 m=1
MP10 GCLK net12 VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MP9 net12 net14 net13 VDD p105 w=0.75u l=0.03u nf=1.0 m=1
MP7 net14 ENL VDD VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MN12 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN11 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 CLKP net3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 ENL net3 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN5 net3 CLKN net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 EN VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN6 net5 ENL VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 net2 SE VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN8 net12 CLKP VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN10 GCLK net12 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN9 net12 net14 VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN7 net14 ENL VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
.ends CGLNPRX8_RVT




.subckt CGLNPSX16_RVT CLK EN GCLK SE VDD VSS
MP15 GCLK net148 VDD VDD p105 w=0.8u l=0.03u nf=1 m=16
MP14 net148 net146 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP2 net1 CLKN net2 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net8 CLKP VDD VDD p105 w=0.7u l=0.03u nf=1 m=1
MP7 ENL net5 net6 VDD p105 w=0.7u l=0.03u nf=1 m=1
MP5 net2 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net146 net9 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP6 net6 SE VDD VDD p105 w=0.7u l=0.03u nf=1 m=1
MP11 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP9 net9 ENL net8 VDD p105 w=0.7u l=0.03u nf=1 m=1
MP12 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP3 net5 net2 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP4 net3 net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MN15 GCLK net148 VSS VSS n105 w=0.42u l=0.03u nf=1 m=16
MN14 net148 net146 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN4 net2 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 ENL SE VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN10 net146 net9 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN7 ENL net5 VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN5 net4 net5 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN8 net9 CLKP VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN11 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN9 net9 ENL VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN2 net1 CLKP net2 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN3 net5 net2 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
.ends CGLNPSX16_RVT




.subckt CGLNPSX2_RVT CLK EN GCLK SE VDD VSS
MN2 net1 CLKP net2 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 net9 ENL VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN11 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN8 net9 CLKP VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN7 ENL net5 VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN6 ENL SE VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN3 net5 net2 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN5 net4 net5 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN10 GCLK net9 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN4 net2 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MP3 net5 net2 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP6 net6 SE VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP5 net2 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net8 CLKP VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP2 net1 CLKN net2 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net3 net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP12 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP9 net9 ENL net8 VDD p105 w=0.6u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP11 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP10 GCLK net9 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP7 ENL net5 net6 VDD p105 w=0.6u l=0.03u nf=1 m=1
.ends CGLNPSX2_RVT




.subckt CGLNPSX4_RVT CLK EN GCLK SE VDD VSS
MP2 net1 CLKN net2 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net8 CLKP VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP7 ENL net5 net6 VDD p105 w=0.6u l=0.03u nf=1 m=1
MP5 net2 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 GCLK net9 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP6 net6 SE VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP11 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP9 net9 ENL net8 VDD p105 w=0.6u l=0.03u nf=1 m=1
MP12 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP3 net5 net2 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP4 net3 net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MN4 net2 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 ENL SE VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN10 GCLK net9 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN7 ENL net5 VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN5 net4 net5 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN8 net9 CLKP VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN11 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN9 net9 ENL VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN2 net1 CLKP net2 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN3 net5 net2 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
.ends CGLNPSX4_RVT




.subckt CGLNPSX8_RVT CLK EN GCLK SE VDD VSS
MP2 net1 CLKN net2 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net8 CLKP VDD VDD p105 w=0.7u l=0.03u nf=1 m=1
MP7 ENL net5 net6 VDD p105 w=0.7u l=0.03u nf=1 m=1
MP5 net2 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 GCLK net9 VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MP6 net6 SE VDD VDD p105 w=0.7u l=0.03u nf=1 m=1
MP11 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP9 net9 ENL net8 VDD p105 w=0.7u l=0.03u nf=1 m=1
MP12 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP3 net5 net2 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP4 net3 net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MN4 net2 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 ENL SE VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN10 GCLK net9 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN7 ENL net5 VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN5 net4 net5 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN8 net9 CLKP VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN11 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN9 net9 ENL VSS VSS n105 w=0.2u l=0.03u nf=1 m=1
MN2 net1 CLKP net2 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN3 net5 net2 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
.ends CGLNPSX8_RVT




.subckt CGLPPRX2_RVT CLK EN GCLK SE VDD VSS
MN8 net7 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net6 ENL net7 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 GCLK net6 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net2 SE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 EN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN11 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN6 net5 ENL VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 net3 CLKP net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 ENL net3 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 CLKN net3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP9 GCLK net6 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP8 net6 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net6 ENL VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 net2 EN net1 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 net1 SE VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP5 net4 ENL VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net3 CLKN net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP4 ENL net3 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP10 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP11 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP3 net2 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends CGLPPRX2_RVT




.subckt CGLPPRX8_RVT CLK EN GCLK SE VDD VSS
MP8 net6 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net3 CLKN net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP4 ENL net3 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP10 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP11 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP3 net2 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net6 ENL VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 net2 EN net1 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 net1 SE VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP9 GCLK net6 VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MP5 net4 ENL VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MN1 net2 SE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 EN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN6 net5 ENL VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 net3 CLKP net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN4 ENL net3 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 CLKN net3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN8 net7 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net6 ENL net7 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 GCLK net6 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
.ends CGLPPRX8_RVT




.subckt CGLPPSX16_RVT CLK EN GCLK SE VDD VSS
MN4 net5 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN10 GCLK net136 VSS VSS n105 w=0.42u l=0.03u nf=1 m=16
MM15 net139 SE VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM13 net136 ENL net137 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 ENL net139 net138 VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 CLKP net5 VSS n105 w=0.3u l=0.03u nf=1 m=1
MM11 net137 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 net138 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN11 CLKP CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 net140 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKN CLKP VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN5 net4 net140 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MM14 net139 SE VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MM12 net136 ENL VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 ENL net139 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 net5 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP2 net1 CLKN net5 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net140 net5 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP4 net3 net140 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 CLKP CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP10 GCLK net136 VDD VDD p105 w=0.8u l=0.03u nf=1 m=16
MP7 ENL net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP12 CLKN CLKP VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MM10 net136 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends CGLPPSX16_RVT




.subckt CGLPPSX2_RVT CLK EN GCLK SE VDD VSS
MM13 net162 ENL net161 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN2 net1 CLKP net5 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN11 CLKP CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN7 ENL net166 net160 VSS n105 w=0.18u l=0.03u nf=1 m=1
MM11 net161 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 net160 net5 VSS VSS n105 w=0.18u l=0.03u nf=1 m=1
MN3 net165 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKN CLKP VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN5 net4 net165 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN10 GCLK net162 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN4 net5 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MM15 net166 SE VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM12 net162 ENL VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net165 net5 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP6 ENL net166 VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP5 net5 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP2 net1 CLKN net5 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net3 net165 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP12 CLKN CLKP VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MM10 net162 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP11 CLKP CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP10 GCLK net162 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP7 ENL net5 VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MM14 net166 SE VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
.ends CGLPPSX2_RVT




.subckt CGLPPSX4_RVT CLK EN GCLK SE VDD VSS
MN5 net4 net140 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN12 CLKN CLKP VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 net140 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN11 CLKP CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN6 net138 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM11 net137 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN2 net1 CLKP net5 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 ENL net139 net138 VSS n105 w=0.4u l=0.03u nf=1 m=1
MM13 net136 ENL net137 VSS n105 w=0.3u l=0.03u nf=1 m=1
MM15 net139 SE VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN4 net5 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN10 GCLK net136 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MM10 net136 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP12 CLKN CLKP VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP4 net3 net140 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net140 net5 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 CLKN net5 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 net5 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 ENL net139 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MM12 net136 ENL VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MM14 net139 SE VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP7 ENL net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 GCLK net136 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP11 CLKP CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends CGLPPSX4_RVT




.subckt CGLPPSX8_RVT CLK EN GCLK SE VDD VSS
MN4 net5 CLKN net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN10 GCLK net136 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MM15 net139 SE VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM13 net136 ENL net137 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 ENL net139 net138 VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 CLKP net5 VSS n105 w=0.3u l=0.03u nf=1 m=1
MM11 net137 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 net138 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN11 CLKP CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 net140 net5 VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN1 net1 EN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN12 CLKN CLKP VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN5 net4 net140 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MM14 net139 SE VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MM12 net136 ENL VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 ENL net139 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 net5 CLKP net3 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP2 net1 CLKN net5 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net140 net5 VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP4 net3 net140 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 CLKP CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP10 GCLK net136 VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MP7 ENL net5 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP12 CLKN CLKP VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP1 net1 EN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MM10 net136 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends CGLPPSX8_RVT




.subckt CLOAD1_RVT A VDD VSS
MN0 VSS A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP0 VDD A VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends CLOAD1_RVT




.subckt DCAP_RVT VDD VSS
MN0 VSS net55 net54 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP0 net55 net54 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
.ends DCAP_RVT



.GLOBAL VDD VSS
.subckt DEC24X1_RVT A0 A1 VDD VSS Y0 Y1 Y2 Y3
MN12 Y1 net438 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN11 Y0 net437 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN8 net423 A0 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN7 net439 net421 net423 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN6 net416 net415 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN10 net428 A0 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN9 net440 A1 net428 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN13 Y2 net439 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 net438 A1 net416 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net409 net415 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net437 net421 net409 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN14 Y3 net440 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net415 A0 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net421 A1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP12 Y1 net438 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP8 net439 net421 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 net440 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP7 net439 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP11 Y0 net437 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP6 net438 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP9 net440 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP13 Y2 net439 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP4 net437 net421 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP3 net437 net415 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 Y3 net440 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP5 net438 net415 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 net421 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net415 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends DEC24X1_RVT



.GLOBAL VDD VSS
.subckt DEC24X2_RVT A0 A1 VDD VSS Y0 Y1 Y2 Y3
MN12 Y1 net438 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 Y0 net437 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN8 net423 A0 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN7 net439 net421 net423 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN6 net416 net415 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN10 net428 A0 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN9 net440 A1 net428 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN13 Y2 net439 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 net438 A1 net416 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net409 net415 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net437 net421 net409 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN14 Y3 net440 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net415 A0 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net421 A1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP12 Y1 net438 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP8 net439 net421 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 net440 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP7 net439 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP11 Y0 net437 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP6 net438 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP9 net440 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP13 Y2 net439 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP4 net437 net421 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP3 net437 net415 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 Y3 net440 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP5 net438 net415 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 net421 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net415 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends DEC24X2_RVT




.subckt DELLN1X2_RVT A VDD VSS Y
MN4 net384 VDD VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN3 net382 VDD net384 VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN1 SA1 A VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MN2 SA2 SA1 net382 VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN8 net398 VDD VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN7 net400 VDD net398 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN5 SA3 SA2 VSS VSS n105 w=0.11u l=0.03u nf=1.0 m=1
MN6 SA4 SA3 net400 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN10 Y SA5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 SA5 SA4 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MP4 net375 VSS VDD VDD p105 w=0.32u l=0.03u nf=1.0 m=1
MP3 net377 VSS net375 VDD p105 w=0.32u l=0.03u nf=1.0 m=1
MP1 SA1 A VDD VDD p105 w=0.23u l=0.03u nf=1.0 m=1
MP2 SA2 SA1 net377 VDD p105 w=0.32u l=0.03u nf=1.0 m=1
MP8 net391 VSS VDD VDD p105 w=0.46u l=0.03u nf=1.0 m=1
MP7 net393 VSS net391 VDD p105 w=0.46u l=0.03u nf=1.0 m=1
MP5 SA3 SA2 VDD VDD p105 w=0.21u l=0.03u nf=1.0 m=1
MP6 SA4 SA3 net393 VDD p105 w=0.46u l=0.03u nf=1.0 m=1
MP10 Y SA5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP9 SA5 SA4 VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
.ends DELLN1X2_RVT




.subckt DELLN2X2_RVT A VDD VSS Y
MN4 net481 VDD VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN3 net480 VDD net481 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MN2 SA2 SA1 net480 VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN8 net471 VDD VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN7 net470 VDD net471 VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN5 SA3 SA2 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MN6 SA4 SA3 net470 VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN12 net463 VDD VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN11 net462 VDD net463 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN9 SA5 SA4 VSS VSS n105 w=0.11u l=0.03u nf=1.0 m=1
MN10 SA6 SA5 net462 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN14 Y SA7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 SA7 SA6 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MP4 net482 VSS VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP3 net483 VSS net482 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 SA1 A VDD VDD p105 w=0.22u l=0.03u nf=1.0 m=1
MP2 SA2 SA1 net483 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net466 VSS VDD VDD p105 w=0.32u l=0.03u nf=1.0 m=1
MP7 net467 VSS net466 VDD p105 w=0.32u l=0.03u nf=1.0 m=1
MP5 SA3 SA2 VDD VDD p105 w=0.23u l=0.03u nf=1.0 m=1
MP6 SA4 SA3 net467 VDD p105 w=0.32u l=0.03u nf=1.0 m=1
MP12 net458 VSS VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP11 net459 VSS net458 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP9 SA5 SA4 VDD VDD p105 w=0.21u l=0.03u nf=1.0 m=1
MP10 SA6 SA5 net459 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP14 Y SA7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 SA7 SA6 VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
.ends DELLN2X2_RVT




.subckt DELLN3X2_RVT A VDD VSS Y
MN4 net638 VDD VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 net640 VDD net638 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN1 SA1 A VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN2 SA2 SA1 net640 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN8 net634 VDD VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN7 net635 VDD net634 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN5 SA3 SA2 VSS VSS n105 w=0.14u l=0.03u nf=1.0 m=1
MN6 SA4 SA3 net635 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 net630 VDD VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN11 net631 VDD net630 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN9 SA5 SA4 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MN10 SA6 SA5 net631 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN16 net626 VDD VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN15 net627 VDD net626 VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN13 SA7 SA6 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MN14 SA8 SA7 net627 VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN20 net622 VDD VSS VSS n105 w=0.23u l=0.03u nf=1.0 m=1
MN19 net623 VDD net622 VSS n105 w=0.23u l=0.03u nf=1.0 m=1
MN17 SA9 SA8 VSS VSS n105 w=0.11u l=0.03u nf=1.0 m=1
MN18 SA10 SA9 net623 VSS n105 w=0.23u l=0.03u nf=1.0 m=1
MN22 Y SA11 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN21 SA11 SA10 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MP4 net617 VSS VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP3 net619 VSS net617 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP1 SA1 A VDD VDD p105 w=0.16u l=0.03u nf=1.0 m=1
MP2 SA2 SA1 net619 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP8 net613 VSS VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP7 net614 VSS net613 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP5 SA3 SA2 VDD VDD p105 w=0.16u l=0.03u nf=1.0 m=1
MP6 SA4 SA3 net614 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP12 net609 VSS VDD VDD p105 w=0.28u l=0.03u nf=1.0 m=1
MP11 net610 VSS net609 VDD p105 w=0.28u l=0.03u nf=1.0 m=1
MP9 SA5 SA4 VDD VDD p105 w=0.14u l=0.03u nf=1.0 m=1
MP10 SA6 SA5 net610 VDD p105 w=0.28u l=0.03u nf=1.0 m=1
MP16 net605 VSS VDD VDD p105 w=0.34u l=0.03u nf=1.0 m=1
MP15 net606 VSS net605 VDD p105 w=0.34u l=0.03u nf=1.0 m=1
MP13 SA7 SA6 VDD VDD p105 w=0.16u l=0.03u nf=1.0 m=1
MP14 SA8 SA7 net606 VDD p105 w=0.34u l=0.03u nf=1.0 m=1
MP20 net601 VSS VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP19 net602 VSS net601 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP17 SA9 SA8 VDD VDD p105 w=0.14u l=0.03u nf=1.0 m=1
MP18 SA10 SA9 net602 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP22 Y SA11 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP21 SA11 SA10 VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
.ends DELLN3X2_RVT




.subckt DFFARX1_RVT CLK D Q QN RSTB VDD VSS
MN8 net294 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net294 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
.ends DFFARX1_RVT




.subckt DFFARX2_RVT CLK D Q QN RSTB VDD VSS
MN8 net294 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net294 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
.ends DFFARX2_RVT




.subckt DFFASRX1_RVT CLK D Q QN RSTB SETB VDD VSS
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 D3 SETB net254 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net253 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN8 net253 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net254 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends DFFASRX1_RVT




.subckt DFFASRX2_RVT CLK D Q QN RSTB SETB VDD VSS
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 D3 SETB net254 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net253 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN8 net253 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net254 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends DFFASRX2_RVT




.subckt DFFASX1_RVT CLK D Q QN SETB VDD VSS
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 D5 D4 VSS VSS n105 w=0.27u l=0.03u nf=1 m=1
MN3 D3 SETB net242 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net242 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP8 D5 D4 VDD VDD p105 w=0.76u l=0.03u nf=1.0 m=1
.ends DFFASX1_RVT




.subckt DFFASX2_RVT CLK D Q QN SETB VDD VSS
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 D5 D4 VSS VSS n105 w=0.27u l=0.03u nf=1 m=1
MN3 D3 SETB net242 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net242 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP8 D5 D4 VDD VDD p105 w=0.76u l=0.03u nf=1.0 m=1
.ends DFFASX2_RVT




.subckt DFFNARX1_RVT CLK D Q QN RSTB VDD VSS
MM19 VDD net7 net211 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net211 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP26 VDD net213 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net213 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net2 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net191 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net7 CLKN net191 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net213 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 net213 CLKP net211 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM18 net211 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net211 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN25 net3 net213 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN23 net213 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net213 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net191 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net7 CLKP net191 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN7 net213 CLKN net211 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends DFFNARX1_RVT




.subckt DFFNARX2_RVT CLK D Q QN RSTB VDD VSS
MM19 VDD net7 net211 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net211 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP26 VDD net213 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net213 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 net191 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net7 CLKN net191 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net213 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 net213 CLKP net211 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM18 net211 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net211 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN25 net3 net213 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN23 net213 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net213 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net191 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net7 CLKP net191 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN7 net213 CLKN net211 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends DFFNARX2_RVT




.subckt DFFNASRNX1_RVT CLK D QN RSTB SETB VDD VSS
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNASRNX1_RVT




.subckt DFFNASRNX2_RVT CLK D QN RSTB SETB VDD VSS
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNASRNX2_RVT




.subckt DFFNASRQX1_RVT CLK D Q RSTB SETB VDD VSS
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNASRQX1_RVT




.subckt DFFNASRQX2_RVT CLK D Q RSTB SETB VDD VSS
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNASRQX2_RVT




.subckt DFFNASRX1_RVT CLK D Q QN RSTB SETB VDD VSS
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNASRX1_RVT




.subckt DFFNASRX2_RVT CLK D Q QN RSTB SETB VDD VSS
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNASRX2_RVT




.subckt DFFNASX1_RVT CLK D Q QN SETB VDD VSS
MM12 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM11 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD net7 net8 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM14 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net8 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends DFFNASX1_RVT




.subckt DFFNASX2_RVT CLK D Q QN SETB VDD VSS
MM12 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM11 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD net7 net8 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM14 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net8 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends DFFNASX2_RVT




.subckt DFFNX1_RVT CLK D Q QN VDD VSS
MN11 net7 net139 net141 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net142 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 net1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN8 net139 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net139 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net141 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net142 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP8 VDD net7 net139 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net139 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP10 net140 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP11 net7 net139 net140 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNX1_RVT




.subckt DFFNX2_RVT CLK D Q QN VDD VSS
MN11 net7 net139 net141 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net142 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 net1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN8 net139 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net139 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 net01 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net141 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net142 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP8 VDD net7 net139 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net139 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 net01 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP10 net140 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP11 net7 net139 net140 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends DFFNX2_RVT




.subckt DFFSSRX1_RVT CLK D Q QN RSTB SETB VDD VSS
MN6 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN01 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 net02 SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN03 net02 D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 IQN net8 net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 net1 CLKN net02 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 IQN CLKP net2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN IQN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN8 net8 IQN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net2 net1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP01 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 net02 RSTB net218 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 net02 D net218 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 net218 SET VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 net226 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP12 IQN net8 net226 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 net1 CLKP net02 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP7 IQN CLKN net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP4 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP14 QN IQN VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP8 net8 IQN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends DFFSSRX1_RVT




.subckt DFFSSRX2_RVT CLK D Q QN RSTB SETB VDD VSS
MN6 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN01 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 net02 SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN03 net02 D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 IQN net8 net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 net1 CLKN net02 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 IQN CLKP net2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN IQN VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN8 net8 IQN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net2 net1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP01 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 net02 RSTB net218 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 net02 D net218 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 net218 SET VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 net226 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP12 IQN net8 net226 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 net1 CLKP net02 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP7 IQN CLKN net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP4 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP14 QN IQN VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP8 net8 IQN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends DFFSSRX2_RVT




.subckt DFFX1_RVT CLK D Q QN VDD VSS
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP12 D5 D4 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 D5 D4 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.30u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.30u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends DFFX1_RVT




.subckt DFFX2_RVT CLK D Q QN VDD VSS
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 D1 D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP12 D5 D4 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN01 D1 D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 D5 D4 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends DFFX2_RVT




.subckt DHFILLH2_RVT VDD VSS
.ends DHFILLH2_RVT




.subckt DHFILLHL2_RVT VDD VSS
.ends DHFILLHL2_RVT




.subckt DHFILLHLHLS11_RVT VDDH VDDL VSS
.ends DHFILLHLHLS11_RVT




.subckt FADDX1_RVT A B CI CO S VDD VSS
MP10 net598 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP12 net607 CI net600 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP11 net600 B net598 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP6 net589 CI VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP7 net589 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP5 net609 B net576 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP8 net589 B VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP4 net576 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP9 net607 net609 net589 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP14 CO net609 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 S net607 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net572 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP3 net609 CI net572 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP2 net572 B VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MN12 net605 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN11 net604 B net605 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN10 net607 CI net604 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN6 net595 CI VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN7 net595 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN5 net579 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN4 net609 B net579 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN13 S net607 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN14 CO net609 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN9 net607 net609 net595 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN3 net573 B VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN1 net573 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN2 net609 CI net573 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN8 net595 B VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
.ends FADDX1_RVT




.subckt FADDX2_RVT A B CI CO S VDD VSS
MP10 net598 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP12 net607 CI net600 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP11 net600 B net598 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP6 net589 CI VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP7 net589 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP5 net609 B net576 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP8 net589 B VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP4 net576 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP9 net607 net609 net589 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP14 CO net609 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP13 S net607 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP1 net572 A VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP3 net609 CI net572 VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MP2 net572 B VDD VDD p105 w=0.62u l=0.03u nf=1.0 m=1
MN12 net605 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN11 net604 B net605 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN10 net607 CI net604 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN6 net595 CI VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN7 net595 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN5 net579 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN4 net609 B net579 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN13 S net607 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN14 CO net609 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN9 net607 net609 net595 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN3 net573 B VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN1 net573 A VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN2 net609 CI net573 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN8 net595 B VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
.ends FADDX2_RVT



.GLOBAL VDD
.subckt FOOT2X16_RVT SLEEP SLEEPOUT VDD VSS VSSG
MP5 SLEEPOUT net71 VDD VDD p105_hvt w=0.8u l=0.03u nf=1 m=16
MP4 net71 SLEEP VDD VDD p105_hvt w=0.8u l=0.03u nf=1.0 m=1
MN10 VSSG net71 VSS VSSG n105_hvt w=0.42u l=0.03u nf=1 m=16
MN3 net71 SLEEP VSSG VSSG n105_hvt w=3.36u l=0.03u nf=8.0 m=1
MN1 SLEEPOUT net71 VSSG VSSG n105_hvt w=0.42u l=0.03u nf=1 m=16
.ends FOOT2X16_RVT



.GLOBAL VDD
.subckt FOOT2X2_RVT SLEEP SLEEPOUT VDD VSS VSSG
MP5 SLEEPOUT net71 VDD VDD p105_hvt w=0.8u l=0.03u nf=1 m=2
MP4 net71 SLEEP VDD VDD p105_hvt w=0.8u l=0.03u nf=1.0 m=1
MN10 VSSG net71 VSS VSSG n105_hvt w=0.42u l=0.03u nf=1 m=2
MN3 net71 SLEEP VSSG VSSG n105_hvt w=0.42u l=0.03u nf=1.0 m=1
MN1 SLEEPOUT net71 VSSG VSSG n105_hvt w=0.42u l=0.03u nf=1 m=2
.ends FOOT2X2_RVT



.GLOBAL VDD
.subckt FOOT2X32_RVT SLEEP SLEEPOUT VDD VSS VSSG
MP5 SLEEPOUT net71 VDD VDD p105_hvt w=0.8u l=0.03u nf=1 m=32
MP4 net71 SLEEP VDD VDD p105_hvt w=0.8u l=0.03u nf=1.0 m=1
MN10 VSSG net71 VSS VSSG n105_hvt w=0.42u l=0.03u nf=1 m=32
MN3 net71 SLEEP VSSG VSSG n105_hvt w=6.72u l=0.03u nf=16.0 m=1
MN1 SLEEPOUT net71 VSSG VSSG n105_hvt w=0.42u l=0.03u nf=1 m=32
.ends FOOT2X32_RVT



.GLOBAL VDD
.subckt FOOT2X4_RVT SLEEP SLEEPOUT VDD VSS VSSG
MP5 SLEEPOUT net71 VDD VDD p105_hvt w=0.8u l=0.03u nf=1 m=4
MP4 net71 SLEEP VDD VDD p105_hvt w=0.8u l=0.03u nf=1.0 m=1
MN10 VSSG net71 VSS VSSG n105_hvt w=0.42u l=0.03u nf=1 m=4
MN3 net71 SLEEP VSSG VSSG n105_hvt w=0.84u l=0.03u nf=2.0 m=1
MN1 SLEEPOUT net71 VSSG VSSG n105_hvt w=0.42u l=0.03u nf=1 m=4
.ends FOOT2X4_RVT



.GLOBAL VDD
.subckt FOOT2X8_RVT SLEEP SLEEPOUT VDD VSS VSSG
MP5 SLEEPOUT net71 VDD VDD p105_hvt w=0.8u l=0.03u nf=1 m=8
MP4 net71 SLEEP VDD VDD p105_hvt w=0.8u l=0.03u nf=1.0 m=1
MN10 VSSG net71 VSS VSSG n105_hvt w=0.42u l=0.03u nf=1.0 m=8
MN3 net71 SLEEP VSSG VSSG n105_hvt w=1.68u l=0.03u nf=4.0 m=1
MN1 SLEEPOUT net71 VSSG VSSG n105_hvt w=0.42u l=0.03u nf=1 m=8
.ends FOOT2X8_RVT




.subckt FOOTX16_RVT SLEEP VDD VSS VSSG
MN8 VSSG SLEEP VSS VSSG n105_hvt w=0.42u l=0.03u nf=1.0 m=16
.ends FOOTX16_RVT




.subckt FOOTX2_RVT SLEEP VDD VSS VSSG
MN8 VSSG SLEEP VSS VSSG n105_hvt w=0.42u l=0.03u nf=1.0 m=2
.ends FOOTX2_RVT




.subckt FOOTX32_RVT SLEEP VDD VSS VSSG
MN8 VSSG SLEEP VSS VSSG n105_hvt w=0.42u l=0.03u nf=1.0 m=32
.ends FOOTX32_RVT




.subckt FOOTX4_RVT SLEEP VDD VSS VSSG
MN8 VSSG SLEEP VSS VSSG n105_hvt w=0.42u l=0.03u nf=1.0 m=4
.ends FOOTX4_RVT




.subckt FOOTX8_RVT SLEEP VDD VSS VSSG
MN8 VSSG SLEEP VSS VSSG n105_hvt w=0.42u l=0.03u nf=1 m=8
.ends FOOTX8_RVT



.GLOBAL VDD
.subckt HADDX1_RVT A0 B0 C1 SO VDD VSS
MP7 C1 net292 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP6 SO net295 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP5 net292 B0 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP4 net292 A0 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP3 net295 net292 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 net295 B0 net288 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net288 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MN6 SO net295 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN7 C1 net292 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 net287 A0 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net292 B0 net287 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net289 net292 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net295 A0 net289 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 net295 B0 net289 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends HADDX1_RVT



.GLOBAL VDD
.subckt HADDX2_RVT A0 B0 C1 SO VDD VSS
MP7 C1 net283 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP6 SO net284 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP5 net283 B0 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP4 net283 A0 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP3 net284 net283 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 net284 B0 net259 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net259 A0 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MN6 SO net284 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN7 C1 net283 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 net282 A0 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net283 B0 net282 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net269 net283 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net284 A0 net269 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 net284 B0 net269 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends HADDX2_RVT




.subckt HEAD2X16_RVT SLEEP SLEEPOUT VDD VDDG VSS
MP1 SLEEPOUT net91 VDDG VDDG p105_lvt w=0.8u l=0.03u nf=1.0 m=16
MP0 net91 SLEEP VDDG VDDG p105_lvt w=0.80u l=0.03u nf=1.0 m=3
MN0 net91 SLEEP VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=3
MN1 SLEEPOUT net91 VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=16
MP2 VDD net91 VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1.0 m=16
.ends HEAD2X16_RVT




.subckt HEAD2X2_RVT SLEEP SLEEPOUT VDD VDDG VSS
MP1 SLEEPOUT net91 VDDG VDDG p105_lvt w=0.8u l=0.03u nf=1.0 m=2
MP0 net91 SLEEP VDDG VDDG p105_lvt w=0.80u l=0.03u nf=1.0 m=1
MN0 net91 SLEEP VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=1
MN1 SLEEPOUT net91 VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=2
MP2 VDD net91 VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1.0 m=2
.ends HEAD2X2_RVT




.subckt HEAD2X32_RVT SLEEP SLEEPOUT VDD VDDG VSS
MP1 SLEEPOUT net91 VDDG VDDG p105_lvt w=0.8u l=0.03u nf=1.0 m=32
MP0 net91 SLEEP VDDG VDDG p105_lvt w=0.80u l=0.03u nf=1.0 m=5
MN0 net91 SLEEP VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=5
MN1 SLEEPOUT net91 VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=32
MP2 VDD net91 VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1.0 m=32
.ends HEAD2X32_RVT




.subckt HEAD2X4_RVT SLEEP SLEEPOUT VDD VDDG VSS
MP1 SLEEPOUT net91 VDDG VDDG p105_lvt w=0.8u l=0.03u nf=1 m=4
MP0 net91 SLEEP VDDG VDDG p105_lvt w=0.80u l=0.03u nf=1.0 m=1
MN0 net91 SLEEP VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=1
MN1 SLEEPOUT net91 VSS VSS n105_lvt w=0.42u l=0.03u nf=1 m=4
MP2 VDD net91 VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1 m=4
.ends HEAD2X4_RVT




.subckt HEAD2X8_RVT SLEEP SLEEPOUT VDD VDDG VSS
MP1 SLEEPOUT net91 VDDG VDDG p105_lvt w=0.8u l=0.03u nf=1.0 m=8
MP0 net91 SLEEP VDDG VDDG p105_lvt w=0.80u l=0.03u nf=1.0 m=2
MN0 net91 SLEEP VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=2
MN1 SLEEPOUT net91 VSS VSS n105_lvt w=0.42u l=0.03u nf=1.0 m=8
MP2 VDD net91 VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1.0 m=8
.ends HEAD2X8_RVT




.subckt HEADX16_RVT SLEEP VDD VDDG VSS
MP0 VDD SLEEP VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1 m=16
.ends HEADX16_RVT




.subckt HEADX2_RVT SLEEP VDD VDDG VSS
MP0 VDD SLEEP VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1.0 m=2
.ends HEADX2_RVT




.subckt HEADX32_RVT SLEEP VDD VDDG VSS
MP0 VDD SLEEP VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1 m=32
.ends HEADX32_RVT




.subckt HEADX4_RVT SLEEP VDD VDDG VSS
MP0 VDD SLEEP VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1 m=4
.ends HEADX4_RVT




.subckt HEADX8_RVT SLEEP VDD VDDG VSS
MP0 VDD SLEEP VDDG VDDG p105_hvt w=0.8u l=0.03u nf=1 m=8
.ends HEADX8_RVT




.subckt IBUFFX16_RVT A VDD VSS Y
MP3 Y 2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=16
MP2 2 1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=3
MP1 1 A VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MN3 Y 2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=16
MN2 2 1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=3
MN1 1 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends IBUFFX16_RVT




.subckt IBUFFX2_RVT A VDD VSS Y
MP3 Y 2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP2 2 1 VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP1 1 A VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MN3 Y 2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN2 2 1 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN1 1 A VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
.ends IBUFFX2_RVT




.subckt IBUFFX32_RVT A VDD VSS Y
MP3 Y 2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=32
MP2 2 1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=6
MP1 1 A VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN3 Y 2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=32
MN2 2 1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=6
MN1 1 A VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
.ends IBUFFX32_RVT




.subckt IBUFFX4_RVT A VDD VSS Y
MP3 Y 2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP2 2 1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 1 A VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MN3 Y 2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN2 2 1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 1 A VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
.ends IBUFFX4_RVT




.subckt IBUFFX8_RVT A VDD VSS Y
MP3 Y net40 VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MP2 net40 net39 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net39 A VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MN3 Y net40 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN2 net40 net39 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net39 A VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends IBUFFX8_RVT




.subckt INVX0_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MN Y A VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends INVX0_RVT




.subckt INVX16_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.8u l=0.03u nf=1 m=16
MN Y A VSS VSS n105 w=0.42u l=0.03u nf=1 m=16
.ends INVX16_RVT




.subckt INVX1_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MN Y A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends INVX1_RVT



.GLOBAL VDD VSS
.subckt INVX2_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN Y A VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
.ends INVX2_RVT




.subckt INVX32_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.8u l=0.03u nf=1 m=32
MN Y A VSS VSS n105 w=0.42u l=0.03u nf=1 m=32
.ends INVX32_RVT




.subckt INVX4_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MN Y A VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
.ends INVX4_RVT




.subckt INVX8_RVT A VDD VSS Y
MP Y A VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MN Y A VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
.ends INVX8_RVT




.subckt ISOLANDAOX1_RVT D ISO Q VDD VDDG VSS
MN1 net77 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 SD net77 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN4 Q ISO1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN3 ISO1 D SD VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MP1 net77 ISO VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 ISO1 net77 VDDG VDDG p105 w=0.18u l=0.03u nf=1.0 m=2
MP3 ISO1 D VDDG VDDG p105 w=0.18u l=0.03u nf=1.0 m=2
MP4 Q ISO1 VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
.ends ISOLANDAOX1_RVT




.subckt ISOLANDAOX2_RVT D ISO Q VDD VDDG VSS
MP3 ISO1 D VDDG VDDG p105 w=0.18u l=0.03u nf=1.0 m=2
MP2 ISO1 net32 VDDG VDDG p105 w=0.18u l=0.03u nf=1.0 m=2
MP1 net32 ISO VDDG VDDG p105 w=0.44u l=0.03u nf=1.0 m=1
MP4 Q ISO1 VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=4
MN1 net32 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 SD net32 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN3 ISO1 D SD VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN4 Q ISO1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=4
.ends ISOLANDAOX2_RVT




.subckt ISOLANDAOX4_RVT D ISO Q VDD VDDG VSS
MP3 ISO1 D VDDG VDDG p105 w=0.18u l=0.03u nf=1.0 m=2
MP2 ISO1 net36 VDDG VDDG p105 w=0.18u l=0.03u nf=1.0 m=2
MP4 Q ISO1 VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=8
MP1 net36 ISO VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=1
MN3 ISO1 D SD VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN4 Q ISO1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=8
MN1 net36 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 SD net36 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
.ends ISOLANDAOX4_RVT




.subckt ISOLANDAOX8_RVT D ISO Q VDD VDDG VSS
MP4 Q ISO1 VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=16
MP3 ISO1 D VDDG VDDG p105 w=0.22u l=0.03u nf=1.0 m=2
MP2 ISO1 net37 VDDG VDDG p105 w=0.22u l=0.03u nf=1.0 m=2
MP1 net37 ISO VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=1
MN2 SD net37 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=2
MN4 Q ISO1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=16
MN1 net37 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 ISO1 D SD VSS n105 w=0.22u l=0.03u nf=1.0 m=2
.ends ISOLANDAOX8_RVT




.subckt ISOLANDX1_RVT D ISO Q VDD VSS
MM25 net101 ISO VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MM22 ISO1 net101 VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MM21 ISO1 D VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MM20 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MM24 net101 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MM23 SD net101 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM19 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM18 ISO1 D SD VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends ISOLANDX1_RVT




.subckt ISOLANDX2_RVT D ISO Q VDD VSS
MM25 net16 ISO VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MM20 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MM21 ISO1 D VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MM22 ISO1 net16 VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MM19 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MM18 ISO1 D SD VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM23 SD net16 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM24 net16 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
.ends ISOLANDX2_RVT




.subckt ISOLANDX4_RVT D ISO Q VDD VSS
MM25 net16 ISO VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MM20 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MM21 ISO1 D VDD VDD p105 w=0.34u l=0.03u nf=1.0 m=1
MM22 ISO1 net16 VDD VDD p105 w=0.34u l=0.03u nf=1.0 m=1
MM23 SD net16 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM18 ISO1 D SD VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM19 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MM24 net16 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
.ends ISOLANDX4_RVT




.subckt ISOLANDX8_RVT D ISO Q VDD VSS
MM25 net16 ISO VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MM20 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=8
MM21 ISO1 D VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MM22 ISO1 net16 VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
MM19 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=8
MM18 ISO1 D SD VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM23 SD net16 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM24 net16 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
.ends ISOLANDX8_RVT




.subckt ISOLORAOX1_RVT D ISO Q VDD VDDG VSS
MN1 net47 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 net46 net47 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN5 Q net54 VSS VSS n105 w=0.21u l=0.03u nf=1 m=2
MN4 net54 ISO VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=2
MN3 net54 net46 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=2
MP1 net47 D VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 net46 net47 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP5 Q net54 VDDG VDDG p105 w=0.40u l=0.03u nf=1 m=2
MP4 net35 ISO VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
MP3 net54 net46 net35 VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
.ends ISOLORAOX1_RVT




.subckt ISOLORAOX2_RVT D ISO Q VDD VDDG VSS
MP3 net32 net34 net33 VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
MP5 Q net32 VDDG VDDG p105 w=0.40u l=0.03u nf=1 m=4
MP4 net33 ISO VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
MP2 net34 net35 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP1 net35 D VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MN3 net32 net34 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=2
MN4 net32 ISO VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=2
MN5 Q net32 VSS VSS n105 w=0.21u l=0.03u nf=1 m=4
MN2 net34 net35 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN1 net35 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
.ends ISOLORAOX2_RVT




.subckt ISOLORAOX4_RVT D ISO Q VDD VDDG VSS
MP2 net32 net33 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP3 net30 net32 net31 VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
MP1 net33 D VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 net31 ISO VDDG VDDG p105 w=0.40u l=0.03u nf=1.0 m=2
MP5 Q net30 VDDG VDDG p105 w=0.40u l=0.03u nf=1 m=8
MN3 net30 net32 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=2
MN2 net32 net33 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN4 net30 ISO VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=2
MN1 net33 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN5 Q net30 VSS VSS n105 w=0.21u l=0.03u nf=1 m=8
.ends ISOLORAOX4_RVT




.subckt ISOLORAOX8_RVT D ISO Q VDD VDDG VSS
MP1 net38 D VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP3 net35 net37 net36 VDDG p105 w=0.42u l=0.03u nf=1.0 m=3
MP2 net37 net38 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP5 Q net35 VDDG VDDG p105 w=0.40u l=0.03u nf=1 m=16
MP4 net36 ISO VDDG VDDG p105 w=0.42u l=0.03u nf=1.0 m=3
MN3 net35 net37 VSS VSS n105 w=0.14u l=0.03u nf=1.0 m=3
MN4 net35 ISO VSS VSS n105 w=0.14u l=0.03u nf=1.0 m=3
MN1 net38 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 net37 net38 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN5 Q net35 VSS VSS n105 w=0.21u l=0.03u nf=1 m=16
.ends ISOLORAOX8_RVT




.subckt ISOLORX1_RVT D ISO Q VDD VSS
MP2 ISO1 D SD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 SD ISO VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MN1 ISO1 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 ISO1 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
.ends ISOLORX1_RVT




.subckt ISOLORX2_RVT D ISO Q VDD VSS
MP2 ISO1 D SD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP1 SD ISO VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MN1 ISO1 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 ISO1 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
.ends ISOLORX2_RVT




.subckt ISOLORX4_RVT D ISO Q VDD VSS
MP2 ISO1 D SD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1 m=4
MP1 SD ISO VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MN2 ISO1 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN1 ISO1 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
.ends ISOLORX4_RVT




.subckt ISOLORX8_RVT D ISO Q VDD VSS
MP2 ISO1 D SD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP3 Q ISO1 VDD VDD p105 w=0.80u l=0.03u nf=1 m=8
MP1 SD ISO VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MN2 ISO1 D VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=2
MN1 ISO1 ISO VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=2
MN3 Q ISO1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
.ends ISOLORX8_RVT




.subckt LARX1_RVT CLK D Q QN RSTB VDD VSS
MP5 net3 IQN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP9 QN net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 Q net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MN5 net3 IQN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 QN net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN10 Q net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
.ends LARX1_RVT




.subckt LARX2_RVT CLK D Q QN RSTB VDD VSS
MP5 net3 IQN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP9 QN net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 Q net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net1 D VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MN5 net3 IQN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 QN net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN10 Q net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
.ends LARX2_RVT




.subckt LASRNX1_RVT CLK D QN RSTB SETB VDD VSS
MN10 net4 IQN VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN11 net3 SETB net4 VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 QN net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MP10 net3 IQN VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP11 net3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.4u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP9 QN net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASRNX1_RVT




.subckt LASRNX2_RVT CLK D QN RSTB SETB VDD VSS
MN10 net4 IQN VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN11 net3 SETB net4 VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 QN net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MP10 net3 IQN VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP11 net3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.4u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP9 QN net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASRNX2_RVT




.subckt LASRQX1_RVT CLK D Q RSTB SETB VDD VSS
MM5 Q net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN10 net4 IQN VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN11 net3 SETB net4 VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MM4 Q net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP10 net3 IQN VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP11 net3 SETB VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASRQX1_RVT




.subckt LASRQX2_RVT CLK D Q RSTB SETB VDD VSS
MM5 Q net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN10 net4 IQN VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN11 net3 SETB net4 VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MM4 Q net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP10 net3 IQN VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP11 net3 SETB VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.6u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASRQX2_RVT




.subckt LASRX1_RVT CLK D Q QN RSTB SETB VDD VSS
MN9 QN net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MM5 Q net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN10 net4 IQN VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN11 net3 SETB net4 VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MP9 QN net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MM4 Q net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP10 net3 IQN VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP11 net3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.4u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASRX1_RVT




.subckt LASRX2_RVT CLK D Q QN RSTB SETB VDD VSS
MN9 QN net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM5 Q net5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN10 net4 IQN VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN11 net3 SETB net4 VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP net1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN7 net5 net3 net6 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN8 net6 RSTB VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net1 RSTB net2 VSS n105 w=0.35u l=0.03u nf=1 m=1
MN4 net5 CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 net2 D VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MP9 QN net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM4 Q net5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP10 net3 IQN VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP11 net3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP8 net5 RSTB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 net5 CLKP IQN VDD p105 w=0.4u l=0.03u nf=1 m=1
MP3 IQN CLKN net1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP2 net1 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MP7 net5 net3 VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 net1 D VDD VDD p105 w=0.52u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASRX2_RVT




.subckt LASX1_RVT CLK D Q QN SETB VDD VSS
MN9 QN FB VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN6 Q FBN VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN10 net4 IQN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN11 FB SETB net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN5 FBN FB VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP D1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN4 FBN CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 D1 D VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MP9 QN FB VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP6 Q FBN VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP10 FB IQN VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 FB SETB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP5 FBN FB VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP4 FBN CLKP IQN VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 IQN CLKN D1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 D1 D VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASX1_RVT




.subckt LASX2_RVT CLK D Q QN SETB VDD VSS
MN9 QN FB VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN6 Q FBN VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN10 net4 IQN VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN11 FB SETB net4 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN5 FBN FB VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 IQN CLKP D1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN4 FBN CLKN IQN VSS n105 w=0.3u l=0.03u nf=1 m=1
MN1 D1 D VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MP9 QN FB VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP6 Q FBN VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP10 FB IQN VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 FB SETB VDD VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP5 FBN FB VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP4 FBN CLKP IQN VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 IQN CLKN D1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP1 D1 D VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LASX2_RVT




.subckt LATCHX1_RVT CLK D Q QN VDD VSS
MN5 TG2 FB1 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MM16 FB1 TG1 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MM14 DN D VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 QN FB1 VSS VSS n105 w='0.42um' l=0.03u nf=1 m=1
MM5 Q TG1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 TG1 CLKP DN VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN4 TG2 CLKN TG1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MP5 TG2 FB1 VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MM17 FB1 TG1 VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MM15 DN D VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP9 QN FB1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MM4 Q TG1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP4 TG2 CLKP TG1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP3 TG1 CLKN DN VDD p105 w=0.4u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LATCHX1_RVT




.subckt LATCHX2_RVT CLK D Q QN VDD VSS
MN5 TG2 FB1 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MM16 FB1 TG1 VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MM14 DN D VSS VSS n105 w=0.3u l=0.03u nf=1 m=1
MN9 QN FB1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM5 Q TG1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN3 TG1 CLKP DN VSS n105 w=0.3u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN4 TG2 CLKN TG1 VSS n105 w=0.3u l=0.03u nf=1 m=1
MP5 TG2 FB1 VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MM17 FB1 TG1 VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MM15 DN D VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP9 QN FB1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM4 Q TG1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP4 TG2 CLKP TG1 VDD p105 w=0.4u l=0.03u nf=1 m=1
MP3 TG1 CLKN DN VDD p105 w=0.4u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
.ends LATCHX2_RVT




.subckt LNANDX1_RVT Q QN RIN SIN VDD VSS
MP3 QN RIN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP4 VDD Q QN VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 Q SIN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 VDD QN Q VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MN3 net161 RIN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 QN Q net161 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 Q QN net151 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net151 SIN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LNANDX1_RVT




.subckt LNANDX2_RVT Q QN RIN SIN VDD VSS
MN1 net10 SIN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN2 Q QN net10 VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN4 QN Q net11 VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN3 net11 RIN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MP2 VDD QN Q VDD p105 w=0.3u l=0.03u nf=1.0 m=2
MP4 VDD Q QN VDD p105 w=0.3u l=0.03u nf=1.0 m=2
MP3 QN RIN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=2
MP1 Q SIN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=2
.ends LNANDX2_RVT




.subckt LSDNENCLSSX1_RVT A EN VDDL VSS Y
MP4 Y net195 net208 VDDL p105 w=0.8u l=0.03u nf=1 m=1
MM10 net208 EN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MP1 net195 A VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MN4 Y net195 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 Y EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net195 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSDNENCLSSX1_RVT




.subckt LSDNENCLSSX2_RVT A EN VDDL VSS Y
MP4 Y net195 net208 VDDL p105 w=0.8u l=0.03u nf=1 m=2
MM10 net208 EN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MP1 net195 A VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MN4 Y net195 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 Y EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net195 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSDNENCLSSX2_RVT




.subckt LSDNENCLSSX4_RVT A EN VDDL VSS Y
MP4 Y net195 net208 VDDL p105 w=0.8u l=0.03u nf=1 m=4
MM10 net208 EN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MP1 net195 A VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MN4 Y net195 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN5 Y EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net195 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSDNENCLSSX4_RVT




.subckt LSDNENCLSSX8_RVT A EN VDDL VSS Y
MP4 Y net195 net208 VDDL p105 w=0.8u l=0.03u nf=1 m=8
MM10 net208 EN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MP1 net195 A VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MN4 Y net195 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN5 Y EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net195 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSDNENCLSSX8_RVT




.subckt LSDNENCLX1_RVT A EN VDDH VDDL VSS Y
MN2 Y net20 VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
MM2 Y EN VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
MN1 net20 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MP3 net46 EN VDDL VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP2 Y net20 net46 VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP1 net20 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
.ends LSDNENCLX1_RVT




.subckt LSDNENCLX2_RVT A EN VDDH VDDL VSS Y
MN3 net61 EN VSS VSS n105 w=0.3u l=0.03u nf=1 m=2
MN5 Y net58 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN2 net61 net57 VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
MN1 net57 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN4 net58 net61 VSS VSS n105 w=0.33u l=0.03u nf=1 m=1
MP5 Y net58 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP4 net58 net61 VDDL VDDL p105 w=0.60u l=0.03u nf=1 m=1
MP3 net59 EN VDDL VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP2 net61 net57 net59 VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP1 net57 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
.ends LSDNENCLX2_RVT




.subckt LSDNENCLX4_RVT A EN VDDH VDDL VSS Y
MP1 net37 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
MP2 net38 net37 net36 VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP3 net36 EN VDDL VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP5 Y net34 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=4
MP4 net34 net38 VDDL VDDL p105 w=0.80u l=0.03u nf=1 m=1
MN1 net37 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN2 net38 net37 VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
MN4 net34 net38 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN3 net38 EN VSS VSS n105 w=0.3u l=0.03u nf=1 m=2
MN5 Y net34 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
.ends LSDNENCLX4_RVT




.subckt LSDNENCLX8_RVT A EN VDDH VDDL VSS Y
MP4 net34 net38 VDDL VDDL p105 w=0.80u l=0.03u nf=1 m=2
MP5 Y net34 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=8
MP3 net36 EN VDDL VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP2 net38 net37 net36 VDDL p105 w=0.75u l=0.03u nf=1.0 m=2
MP1 net37 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
MN3 net38 EN VSS VSS n105 w=0.35u l=0.03u nf=1 m=2
MN4 net34 net38 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 Y net34 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN1 net37 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN2 net38 net37 VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
.ends LSDNENCLX8_RVT




.subckt LSDNENSSX1_RVT A EN VDDL VSS Y
MM10 net167 EN VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP4 Y SA3 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA3 SA2 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA2 SA1 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 SA1 A VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP5 Y net167 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MM11 net167 EN VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN4 Y SA3 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA3 SA2 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA2 SA1 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 VSSV net167 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN1 SA1 A VSSV VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends LSDNENSSX1_RVT




.subckt LSDNENSSX2_RVT A EN VDDL VSS Y
MM10 net167 EN VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP4 Y SA3 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP3 SA3 SA2 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA2 SA1 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 SA1 A VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP5 Y net167 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MM11 net167 EN VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN4 Y SA3 VSSV VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 SA3 SA2 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA2 SA1 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 VSSV net167 VSS VSS n105 w=0.42u l=0.03u nf=1 m=6
MN1 SA1 A VSSV VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends LSDNENSSX2_RVT




.subckt LSDNENSSX4_RVT A EN VDDL VSS Y
MM10 net167 EN VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP4 Y SA3 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=4
MP3 SA3 SA2 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA2 SA1 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 SA1 A VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP5 Y net167 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=4
MM11 net167 EN VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN4 Y SA3 VSSV VSS n105 w=0.42u l=0.03u nf=1 m=4
MN3 SA3 SA2 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA2 SA1 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 VSSV net167 VSS VSS n105 w=0.42u l=0.03u nf=1 m=6
MN1 SA1 A VSSV VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends LSDNENSSX4_RVT




.subckt LSDNENSSX8_RVT A EN VDDL VSS Y
MM10 net167 EN VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP4 Y SA3 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=8
MP3 SA3 SA2 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP2 SA2 SA1 VDDL VDDL p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 SA1 A VDDL VDDL p105 w=0.52u l=0.03u nf=1.0 m=1
MP5 Y net167 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=6
MM11 net167 EN VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN4 Y SA3 VSSV VSS n105 w=0.42u l=0.03u nf=1 m=8
MN3 SA3 SA2 VSSV VSS n105 w=0.42u l=0.03u nf=1 m=2
MN2 SA2 SA1 VSSV VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 VSSV net167 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN1 SA1 A VSSV VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends LSDNENSSX8_RVT




.subckt LSDNENX1_RVT A EN VDDH VDDL VSS Y
MN0 net31 EN VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN2 Y net20 net21 VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN3 net21 net31 VSS VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN1 net20 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MP0 net31 EN VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=1
MP3 Y net31 VDDL VDDL p105 w=0.66u l=0.03u nf=1.0 m=1
MP2 Y net20 VDDL VDDL p105 w=0.66u l=0.03u nf=1.0 m=1
MP1 net20 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
.ends LSDNENX1_RVT




.subckt LSDNENX2_RVT A EN VDDH VDDL VSS Y
MN0 net31 EN VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN5 Y net24 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN2 net35 net20 net21 VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN3 net21 net31 VSS VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN1 net20 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN4 net24 net35 VSS VSS n105 w=0.33u l=0.03u nf=1 m=1
MP0 net31 EN VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=1
MP5 Y net24 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP4 net24 net35 VDDL VDDL p105 w=0.60u l=0.03u nf=1 m=1
MP3 net35 net31 VDDL VDDL p105 w=0.66u l=0.03u nf=1.0 m=1
MP2 net35 net20 VDDL VDDL p105 w=0.66u l=0.03u nf=1.0 m=1
MP1 net20 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
.ends LSDNENX2_RVT




.subckt LSDNENX4_RVT A EN VDDH VDDL VSS Y
MN0 net31 EN VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN5 Y net24 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN2 net35 net20 net21 VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN3 net21 net31 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN1 net20 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN4 net24 net35 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MP0 net31 EN VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=1
MP5 Y net24 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=4
MP4 net24 net35 VDDL VDDL p105 w=0.80u l=0.03u nf=1 m=1
MP3 net35 net31 VDDL VDDL p105 w=0.7u l=0.03u nf=1.0 m=1
MP2 net35 net20 VDDL VDDL p105 w=0.66u l=0.03u nf=1.0 m=1
MP1 net20 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
.ends LSDNENX4_RVT




.subckt LSDNENX8_RVT A EN VDDH VDDL VSS Y
MN0 net31 EN VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN5 Y net24 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN2 net39 net20 net21 VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN3 net21 net31 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN1 net20 A VSS VSS n105 w=0.17u l=0.03u nf=1.0 m=1
MN4 net24 net39 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MP0 net31 EN VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=1
MP5 Y net24 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=8
MP4 net24 net39 VDDL VDDL p105 w=0.80u l=0.03u nf=1 m=2
MP3 net39 net31 VDDL VDDL p105 w=0.7u l=0.03u nf=1.0 m=1
MP2 net39 net20 VDDL VDDL p105 w=0.66u l=0.03u nf=1.0 m=1
MP1 net20 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=2
.ends LSDNENX8_RVT



.GLOBAL VSS
.subckt LSDNSSX1_RVT A VDDL VSS Y
MP2 Y AN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=1
MP1 AN A VDDL VDDL p105 w=0.3u l=0.03u nf=1 m=1
MN2 Y AN VSS VSS n105 w=0.26u l=0.03u nf=1 m=1
MN1 AN A VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
.ends LSDNSSX1_RVT



.GLOBAL VSS
.subckt LSDNSSX2_RVT A VDDL VSS Y
MP2 Y AN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP1 AN A VDDL VDDL p105 w=0.65u l=0.03u nf=1.0 m=1
MN2 Y AN VSS VSS n105 w=0.26u l=0.03u nf=1 m=2
MN1 AN A VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
.ends LSDNSSX2_RVT



.GLOBAL VSS
.subckt LSDNSSX4_RVT A VDDL VSS Y
MP2 Y AN VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=4
MP1 AN A VDDL VDDL p105 w=0.8u l=0.03u nf=1.0 m=1
MN2 Y AN VSS VSS n105 w=0.26u l=0.03u nf=1 m=4
MN1 AN A VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
.ends LSDNSSX4_RVT




.subckt LSDNSSX8_RVT A VDDL VSS Y
MP2 Y AN VDDL VDD p105 w=0.8u l=0.03u nf=1 m=8
MP1 AN A VDDL VDD p105 w=0.8u l=0.03u nf=1 m=4
MN2 Y AN VSS VSS n105 w=0.26u l=0.03u nf=1 m=8
MN1 AN A VSS VSS n105 w=0.26u l=0.03u nf=1 m=4
.ends LSDNSSX8_RVT




.subckt LSDNX1_RVT A VDDH VDDL VSS Y
MM3 net85 net84 VSS VSS n105 w=0.37u l=0.03u nf=1.0 m=1
MM4 Y net85 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM2 net84 net82 VSS VSS n105 w=0.1u l=0.03u nf=1 m=1
MM1 net82 A VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MP4 Y net85 VDDL VDDL p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net85 net84 VDDL VDDL p105 w=0.5u l=0.03u nf=1.0 m=1
MP1 net82 A VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP2 net84 net82 VDDL VDDL p105 w=0.6u l=0.03u nf=1.0 m=1
.ends LSDNX1_RVT




.subckt LSDNX2_RVT A VDDH VDDL VSS Y
MM3 net85 net84 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM4 Y net85 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM2 net84 net82 VSS VSS n105 w=0.1u l=0.03u nf=1 m=1
MM1 net82 A VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MP4 Y net85 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP3 net85 net84 VDDL VDDL p105 w=0.5u l=0.03u nf=1.0 m=1
MP1 net82 A VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP2 net84 net82 VDDL VDDL p105 w=0.3u l=0.03u nf=1.0 m=1
.ends LSDNX2_RVT




.subckt LSDNX4_RVT A VDDH VDDL VSS Y
MM3 net85 net84 VSS VSS n105 w=0.5u l=0.03u nf=1.0 m=1
MM4 Y net85 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MM2 net84 net82 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MM1 net82 A VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MP4 Y net85 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=4
MP3 net85 net84 VDDL VDDL p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net82 A VDDH VDDH p105 w=0.35u l=0.03u nf=1.0 m=1
MP2 net84 net82 VDDL VDDL p105 w=0.6u l=0.03u nf=1.0 m=1
.ends LSDNX4_RVT




.subckt LSDNX8_RVT A VDDH VDDL VSS Y
MM3 net85 net84 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM4 Y net85 VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MM2 net84 net82 VSS VSS n105 w=0.12u l=0.03u nf=1.0 m=1
MM1 net82 A VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MP4 Y net85 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=8
MP3 net85 net84 VDDL VDDL p105 w=0.8u l=0.03u nf=1 m=2
MP1 net82 A VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP2 net84 net82 VDDL VDDL p105 w=0.5u l=0.03u nf=1.0 m=1
.ends LSDNX8_RVT




.subckt LSUPENCLX1_RVT A EN VDDH VDDL VSS Y
MP4 net79 EN VDDH VDDH p105 w=0.42u l=0.03u nf=1.0 m=1
MP6 net46 A VDDL VDDL p105 w=0.40u l=0.03u nf=1.0 m=2
MP3 Y net69 net79 VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net76 net69 net79 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP2 net69 net76 net79 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MN4 Y EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net76 net46 VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN6 net46 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN3 Y net69 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 net69 A VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
.ends LSUPENCLX1_RVT




.subckt LSUPENCLX2_RVT A EN VDDH VDDL VSS Y
MP4 net79 EN VDDH VDDH p105 w=0.27u l=0.03u nf=1.0 m=2
MP6 net46 A VDDL VDDL p105 w=0.40u l=0.03u nf=1.0 m=2
MP3 Y net69 net79 VDDH p105 w=0.8u l=0.03u nf=1.0 m=2
MP1 net76 net69 net79 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP2 net69 net76 net79 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MN4 Y EN VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=2
MN1 net76 net46 VSS VSS n105 w=0.41u l=0.03u nf=1.0 m=1
MN6 net46 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN3 Y net69 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN2 net69 A VSS VSS n105 w=0.41u l=0.03u nf=1.0 m=1
.ends LSUPENCLX2_RVT




.subckt LSUPENCLX4_RVT A EN VDDH VDDL VSS Y
MP4 net122 EN VDDH VDDH p105 w=0.40u l=0.03u nf=1.0 m=2
MP6 net129 net116 net122 VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net128 A VDDL VDDL p105 w=0.28u l=0.03u nf=1.0 m=1
MP5 net116 net124 net122 VDDH p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 net126 net124 net122 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP3 net124 net126 net122 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP7 Y net129 net122 VDDH p105 w=0.8u l=0.03u nf=1.0 m=4
MN4 Y EN VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=2
MN2 net126 net128 VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN1 net128 A VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN5 net116 net124 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN3 net124 A VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN7 Y net129 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN6 net129 net116 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSUPENCLX4_RVT




.subckt LSUPENCLX8_RVT A EN VDDH VDDL VSS Y
MP2 net90 net89 net86 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP7 Y net87 net86 VDDH p105 w=0.8u l=0.03u nf=1.0 m=8
MP3 net89 net90 net86 VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP5 net88 net89 net86 VDDH p105 w=0.60u l=0.03u nf=1.0 m=1
MP6 net87 net88 net86 VDDH p105 w=0.8u l=0.03u nf=1.0 m=2
MP4 net86 EN VDDH VDDH p105 w=0.80u l=0.03u nf=1.0 m=8
MP1 net91 A VDDL VDDL p105 w=0.40u l=0.03u nf=1.0 m=2
MN6 net87 net88 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN7 Y net87 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=8
MN4 Y EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=8
MN3 net89 A VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN2 net90 net91 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 net88 net89 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN1 net91 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
.ends LSUPENCLX8_RVT




.subckt LSUPENX1_RVT A EN VDDH VDDL VSS Y
MP1 net26 EN VDDH VDDH p105 w=0.7u l=0.03u nf=1.0 m=1
MP5 Y net26 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net21 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP6 Y net29 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net16 net29 VDDH VDDH p105 w=0.21u l=0.03u nf=1.0 m=1
MP4 net29 net16 VDDH VDDH p105 w=0.21u l=0.03u nf=1.0 m=1
MN1 net26 EN VSS VSS n105 w=0.1u l=0.03u nf=1.0 m=1
MN5 net28 net26 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN3 net16 net21 net28 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 net21 A net28 VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN6 Y net29 net28 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 net29 A net28 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSUPENX1_RVT




.subckt LSUPENX2_RVT A EN VDDH VDDL VSS Y
MP7 net31 net38 VDDH VDDH p105 w=0.8u l=0.03u nf=1 m=1
MP1 net34 EN VDDH VDDH p105 w=0.7u l=0.03u nf=1.0 m=1
MP6 net38 net39 VDDH VDDH p105 w=0.1u l=0.03u nf=1 m=1
MP5 Y net34 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=2
MP2 net37 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP8 Y net31 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=2
MP3 net35 net39 VDDH VDDH p105 w=0.18u l=0.03u nf=1.0 m=1
MP4 net39 net35 VDDH VDDH p105 w=0.18u l=0.03u nf=1.0 m=1
MN7 net31 net38 net33 VSS n105 w=0.3u l=0.03u nf=1 m=1
MN6 net38 net39 net33 VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net34 EN VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN5 net33 net34 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN3 net35 net37 net33 VSS n105 w=0.56u l=0.03u nf=1.0 m=1
MN2 net37 A net33 VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN8 Y net31 net33 VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN4 net39 A net33 VSS n105 w=0.56u l=0.03u nf=1.0 m=1
.ends LSUPENX2_RVT




.subckt LSUPENX4_RVT A EN VDDH VDDL VSS Y
MP7 net35 net36 VDDH VDDH p105 w=0.8u l=0.03u nf=1 m=1
MP1 net30 EN VDDH VDDH p105 w=0.7u l=0.03u nf=1.0 m=1
MP6 net36 net33 VDDH VDDH p105 w=0.2u l=0.03u nf=1 m=1
MP5 Y net30 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=4
MP2 net28 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP8 Y net35 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=4
MP3 net22 net33 VDDH VDDH p105 w=0.18u l=0.03u nf=1.0 m=1
MP4 net33 net22 VDDH VDDH p105 w=0.18u l=0.03u nf=1.0 m=1
MN7 net35 net36 net37 VSS n105 w=0.42u l=0.03u nf=1 m=1
MN6 net36 net33 net37 VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net30 EN VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN5 net37 net30 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN3 net22 net28 net37 VSS n105 w=0.45u l=0.03u nf=1.0 m=1
MN2 net28 A net37 VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN8 Y net35 net37 VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN4 net33 A net37 VSS n105 w=0.45u l=0.03u nf=1.0 m=1
.ends LSUPENX4_RVT




.subckt LSUPENX8_RVT A EN VDDH VDDL VSS Y
MP7 net45 net46 VDDH VDDH p105 w=0.8u l=0.03u nf=1 m=2
MP1 net40 EN VDDH VDDH p105 w=0.7u l=0.03u nf=1.0 m=1
MP6 net46 net43 VDDH VDDH p105 w=0.2u l=0.03u nf=1 m=1
MP5 Y net40 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=8
MP2 net38 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP8 Y net45 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=8
MP3 net31 net43 VDDH VDDH p105 w=0.18u l=0.03u nf=1.0 m=1
MP4 net43 net31 VDDH VDDH p105 w=0.18u l=0.03u nf=1.0 m=1
MN7 net45 net46 net47 VSS n105 w=0.42u l=0.03u nf=1 m=2
MN6 net46 net43 net47 VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net40 EN VSS VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN5 net47 net40 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=8
MN3 net31 net38 net47 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 net38 A net47 VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN8 Y net45 net47 VSS n105 w=0.42u l=0.03u nf=1.0 m=8
MN4 net43 A net47 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends LSUPENX8_RVT




.subckt LSUPX1_RVT A VDDH VDDL VSS Y
MP1 net13 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP4 Y net16 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net14 net16 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP3 net16 net14 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MN2 net14 net13 VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN1 net13 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN4 Y net16 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net16 A VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
.ends LSUPX1_RVT




.subckt LSUPX2_RVT A VDDH VDDL VSS Y
MP6 Y net52 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=2
MP5 net52 net51 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net41 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP4 net51 net44 VDDH VDDH p105 w=0.21u l=0.03u nf=1.0 m=1
MP2 net53 net44 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP3 net44 net53 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MN6 Y net52 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN5 net52 net51 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net53 net41 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN1 net41 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN4 net51 net44 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net44 A VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
.ends LSUPX2_RVT




.subckt LSUPX4_RVT A VDDH VDDL VSS Y
MP6 Y net1 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=4
MP5 net1 net2 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net5 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP4 net2 net3 VDDH VDDH p105 w=0.2u l=0.03u nf=1.0 m=1
MP2 net4 net3 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP3 net3 net4 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MN6 Y net1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN5 net1 net2 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net4 net5 VSS VSS n105 w=0.48u l=0.03u nf=1.0 m=1
MN1 net5 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN4 net2 net3 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net3 A VSS VSS n105 w=0.48u l=0.03u nf=1.0 m=1
.ends LSUPX4_RVT




.subckt LSUPX8_RVT A VDDH VDDL VSS Y
MP3 net60 net61 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP2 net61 net60 VDDH VDDH p105 w=0.28u l=0.03u nf=1.0 m=1
MP4 net59 net60 VDDH VDDH p105 w=0.2u l=0.03u nf=1.0 m=1
MP1 net62 A VDDL VDDL p105 w=0.4u l=0.03u nf=1.0 m=2
MP5 net58 net59 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=2
MP6 Y net58 VDDH VDDH p105 w=0.8u l=0.03u nf=1.0 m=8
MN3 net60 A VSS VSS n105 w=0.48u l=0.03u nf=1.0 m=1
MN4 net59 net60 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net62 A VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=2
MN2 net61 net62 VSS VSS n105 w=0.48u l=0.03u nf=1.0 m=1
MN5 net58 net59 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=2
MN6 Y net58 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=8
.ends LSUPX8_RVT




.subckt MUX21X1_RVT A1 A2 S0 VDD VSS Y
MP1 net1 S0 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP3 net3 A1 net2 VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP6 Y net3 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net2 S0 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP5 net3 A2 net5 VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP4 net5 net1 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MN3 net4 net1 VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN2 net3 A1 net4 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN1 net1 S0 VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN6 Y net3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 net6 S0 VSS VSS n105 w=0.24u l=0.03u nf=1.0 m=1
MN4 net3 A2 net6 VSS n105 w=0.24u l=0.03u nf=1.0 m=1
.ends MUX21X1_RVT




.subckt MUX21X2_RVT A1 A2 S0 VDD VSS Y
MP1 net1 S0 VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP3 net3 A1 net2 VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP6 Y net3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP2 net2 S0 VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP5 net3 A2 net5 VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP4 net5 net1 VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MN3 net4 net1 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN2 net3 A1 net4 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN1 net1 S0 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN6 Y net3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN5 net6 S0 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN4 net3 A2 net6 VSS n105 w=0.28u l=0.03u nf=1.0 m=1
.ends MUX21X2_RVT




.subckt MUX41X1_RVT A1 A2 A3 A4 S0 S1 VDD VSS Y
MN9 Y yn VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MNT2 A3A4 S0 yn VSS n105 w=0.30u l=0.03u nf=1 m=1
MNT1 A1A2 NS0 yn VSS n105 w=0.30u l=0.03u nf=1 m=1
MNS0 NS0 S0 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN7 8 A4 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 A3A4 S1 8 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 6 A3 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN6 A3A4 NS1 6 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 4 A2 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN3 A1A2 S1 4 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 2 A1 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 A1A2 NS1 2 VSS n105 w=0.30u l=0.03u nf=1 m=1
MNS1 NS1 S1 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP9 Y yn VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MPT2 A3A4 NS0 yn VDD p105 w=0.50u l=0.03u nf=1 m=1
MPT1 A1A2 S0 yn VDD p105 w=0.50u l=0.03u nf=1 m=1
MPS0 NS0 S0 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP7 7 A4 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP8 A3A4 NS1 7 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP5 5 A3 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP6 A3A4 S1 5 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP4 A1A2 NS1 3 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP3 3 A2 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP2 A1A2 S1 1 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP1 1 A1 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MPS1 NS1 S1 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
.ends MUX41X1_RVT




.subckt MUX41X2_RVT A1 A2 A3 A4 S0 S1 VDD VSS Y
MN9 Y yn VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MNT2 A3A4 S0 yn VSS n105 w=0.38u l=0.03u nf=1 m=1
MNT1 A1A2 NS0 yn VSS n105 w=0.38u l=0.03u nf=1 m=1
MNS0 NS0 S0 VSS VSS n105 w=0.38u l=0.03u nf=1 m=1
MN7 8 A4 VSS VSS n105 w=0.38u l=0.03u nf=1 m=1
MN8 A3A4 S1 8 VSS n105 w=0.38u l=0.03u nf=1 m=1
MN5 6 A3 VSS VSS n105 w=0.38u l=0.03u nf=1 m=1
MN6 A3A4 NS1 6 VSS n105 w=0.38u l=0.03u nf=1 m=1
MN4 4 A2 VSS VSS n105 w=0.38u l=0.03u nf=1 m=1
MN3 A1A2 S1 4 VSS n105 w=0.38u l=0.03u nf=1 m=1
MN1 2 A1 VSS VSS n105 w=0.38u l=0.03u nf=1 m=1
MN2 A1A2 NS1 2 VSS n105 w=0.38u l=0.03u nf=1 m=1
MNS1 NS1 S1 VSS VSS n105 w=0.38u l=0.03u nf=1 m=1
MP9 Y yn VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MPT2 A3A4 NS0 yn VDD p105 w=0.50u l=0.03u nf=1 m=1
MPT1 A1A2 S0 yn VDD p105 w=0.50u l=0.03u nf=1 m=1
MPS0 NS0 S0 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP7 7 A4 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP8 A3A4 NS1 7 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP5 5 A3 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP6 A3A4 S1 5 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP4 A1A2 NS1 3 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP3 3 A2 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MP2 A1A2 S1 1 VDD p105 w=0.50u l=0.03u nf=1 m=1
MP1 1 A1 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
MPS1 NS1 S1 VDD VDD p105 w=0.50u l=0.03u nf=1 m=1
.ends MUX41X2_RVT




.subckt NAND2X0_RVT A1 A2 VDD VSS Y
MN1 Y A1 SA1 VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MP2 Y A2 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 Y A1 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends NAND2X0_RVT




.subckt NAND2X1_RVT A1 A2 VDD VSS Y
MN2 SA1 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 Y2 Y1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP4 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 Y2 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
.ends NAND2X1_RVT




.subckt NAND2X2_RVT A1 A2 VDD VSS Y
MN2 SA1 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN3 Y2 Y1 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP4 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP3 Y2 Y1 VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
.ends NAND2X2_RVT




.subckt NAND2X4_RVT A1 A2 VDD VSS Y
MN2 SA1 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN3 Y2 Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP4 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MP3 Y2 Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NAND2X4_RVT




.subckt NAND3X0_RVT A1 A2 A3 VDD VSS Y
MP3 Y A3 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP2 Y A2 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP1 Y A1 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.40u l=0.03u nf=1.0 m=1
MN3 SA2 A3 VSS VSS n105 w=0.40u l=0.03u nf=1.0 m=1
MN1 Y A1 SA1 VSS n105 w=0.40u l=0.03u nf=1.0 m=1
.ends NAND3X0_RVT




.subckt NAND3X1_RVT A1 A2 A3 VDD VSS Y
MN4 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM17 Y2 Y1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA2 A3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP4 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MM16 Y2 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.25u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.25u l=0.03u nf=1.0 m=1
MP3 Y1 A3 VDD VDD p105 w=0.25u l=0.03u nf=1.0 m=1
.ends NAND3X1_RVT




.subckt NAND3X2_RVT A1 A2 A3 VDD VSS Y
MP4 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MM16 Y2 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP3 Y1 A3 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MM17 Y2 Y1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN3 SA2 A3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends NAND3X2_RVT




.subckt NAND3X4_RVT A1 A2 A3 VDD VSS Y
MN4 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MM17 Y2 Y1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN3 SA2 A3 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP3 Y1 A3 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP4 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MP2 Y1 A2 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MM16 Y2 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
.ends NAND3X4_RVT




.subckt NAND4X0_RVT A1 A2 A3 A4 VDD VSS Y
MP3 Y A3 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 Y A2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP1 Y A1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 Y A4 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MN1 Y A1 SA1 VSS n105 w=0.52u l=0.03u nf=1.0 m=1
MN3 SA2 A3 SA3 VSS n105 w=0.52u l=0.03u nf=1.0 m=1
MN4 SA3 A4 VSS VSS n105 w=0.52u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.52u l=0.03u nf=1.0 m=1
.ends NAND4X0_RVT




.subckt NAND4X1_RVT A1 A2 A3 A4 VDD VSS Y
MM2 Y net15 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP4 Y1 A4 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP1 Y1 A1 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP5 net15 Y1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP3 Y1 A3 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP2 Y1 A2 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MM1 Y net15 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN4 SA3 A4 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA2 A3 SA3 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 net15 Y1 VSS VSS n105 w=0.20u l=0.03u nf=1 m=1
MN1 Y1 A1 SA1 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 SA1 A2 SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends NAND4X1_RVT




.subckt NBUFFX16_RVT A VDD VSS Y
MP2 Y AN VDD VDD p105 w=0.8u l=0.03u nf=1 m=16
MP1 AN A VDD VDD p105 w=0.8u l=0.03u nf=1 m=3
MN2 Y AN VSS VSS n105 w=0.42u l=0.03u nf=1 m=16
MN1 AN A VSS VSS n105 w=0.42u l=0.03u nf=1 m=3
.ends NBUFFX16_RVT




.subckt NBUFFX2_RVT A VDD VSS Y
MP2 Y AN VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP1 AN A VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MN2 Y AN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN1 AN A VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
.ends NBUFFX2_RVT




.subckt NBUFFX32_RVT A VDD VSS Y
MP2 Y AN VDD VDD p105 w=0.8u l=0.03u nf=1 m=32
MP1 AN A VDD VDD p105 w=0.8u l=0.03u nf=1 m=5
MN2 Y AN VSS VSS n105 w=0.42u l=0.03u nf=1 m=32
MN1 AN A VSS VSS n105 w=0.42u l=0.03u nf=1 m=5
.ends NBUFFX32_RVT




.subckt NBUFFX4_RVT A VDD VSS Y
MP2 Y AN VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP1 AN A VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MN2 Y AN VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN1 AN A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends NBUFFX4_RVT




.subckt NBUFFX8_RVT A VDD VSS Y
MP2 Y AN VDD VDD p105 w=0.8u l=0.03u nf=1 m=8
MP1 AN A VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN2 Y AN VSS VSS n105 w=0.42u l=0.03u nf=1 m=8
MN1 AN A VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
.ends NBUFFX8_RVT



.GLOBAL VSS
.subckt NMT1_RVT D G S VDD VSS
MN0 D G S VSS n105 w=0.42u l=0.03u nf=1.0 m=1
.ends NMT1_RVT



.GLOBAL VSS
.subckt NMT2_RVT D G S VDD VSS
MN0 D G S VSS n105 w=0.42u l=0.03u nf=1 m=2
.ends NMT2_RVT



.GLOBAL VSS
.subckt NMT3_RVT D G S VDD VSS
MN0 D G S VSS n105 w=0.42u l=0.03u nf=1 m=4
.ends NMT3_RVT




.subckt NOR2X0_RVT A1 A2 VDD VSS Y
MN4 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MP4 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net84 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net84 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR2X0_RVT




.subckt NOR2X1_RVT A1 A2 VDD VSS Y
MN4 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MP4 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net84 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net84 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR2X1_RVT




.subckt NOR2X2_RVT A1 A2 VDD VSS Y
MN4 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN3 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MP4 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP3 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net84 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net84 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR2X2_RVT




.subckt NOR2X4_RVT A1 A2 VDD VSS Y
MN4 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN3 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MP4 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MP3 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net84 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net84 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR2X4_RVT




.subckt NOR3X0_RVT A1 A2 A3 VDD VSS Y
MN5 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MP5 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP4 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net93 A2 net94 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 net94 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA1 A3 net93 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR3X0_RVT




.subckt NOR3X1_RVT A1 A2 A3 VDD VSS Y
MN5 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN4 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MP5 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP4 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net93 A2 net94 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 net94 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA1 A3 net93 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR3X1_RVT




.subckt NOR3X2_RVT A1 A2 A3 VDD VSS Y
MN5 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN4 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MP5 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP4 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net93 A2 net94 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 net94 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA1 A3 net93 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR3X2_RVT




.subckt NOR3X4_RVT A1 A2 A3 VDD VSS Y
MN5 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=4
MN4 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.14u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.14u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.14u l=0.03u nf=1.0 m=1
MP5 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=4
MP4 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net93 A2 net94 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 net94 A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP3 SA1 A3 net93 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends NOR3X4_RVT




.subckt NOR4X0_RVT A1 A2 A3 A4 VDD VSS Y
MN6 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN4 SA1 A4 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MP6 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP5 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net135 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net138 A3 net137 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net137 A2 net135 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP4 SA1 A4 net138 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends NOR4X0_RVT




.subckt NOR4X1_RVT A1 A2 A3 A4 VDD VSS Y
MN6 Y SA2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN5 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 SA1 A1 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN4 SA1 A4 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MP6 Y SA2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP5 SA2 SA1 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net135 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net138 A3 net137 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net137 A2 net135 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP4 SA1 A4 net138 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends NOR4X1_RVT




.subckt OA21X1_RVT A1 A2 A3 VDD VSS Y
MP3 net6 A3 VDD VDD p105 w=0.25u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP7 Y net6 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MN7 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net6 A3 net2 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
.ends OA21X1_RVT




.subckt OA21X2_RVT A1 A2 A3 VDD VSS Y
MP3 net7 A3 VDD VDD p105 w=0.24u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP2 net7 A2 net1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN3 net7 A3 net2 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
.ends OA21X2_RVT




.subckt OA221X1_RVT A1 A2 A3 A4 A5 VDD VSS Y
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.41u l=0.03u nf=1.0 m=1
MP7 Y net6 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.41u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.41u l=0.03u nf=1.0 m=1
MP5 net6 A5 VDD VDD p105 w=0.23u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.41u l=0.03u nf=1.0 m=1
.ends OA221X1_RVT




.subckt OA221X2_RVT A1 A2 A3 A4 A5 VDD VSS Y
MP2 net6 A2 net1 VDD p105 w=0.44u l=0.03u nf=1.0 m=1
MP5 net6 A5 VDD VDD p105 w=0.23u l=0.03u nf=1.0 m=1
MP7 Y net6 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP4 net6 A4 net3 VDD p105 w=0.44u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.44u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.44u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN7 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN5 net6 A5 net4 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN4 net4 A4 net2 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN3 net4 A3 net2 VSS n105 w=0.36u l=0.03u nf=1.0 m=1
.ends OA221X2_RVT




.subckt OA222X1_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MP1 net1 A1 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP5 net5 A5 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP7 Y net6 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP6 net6 A6 net5 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 net6 A6 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
.ends OA222X1_RVT




.subckt OA222X2_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MP4 net6 A4 net3 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP5 net5 A5 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP6 net6 A6 net5 VDD p105 w=0.42u l=0.03u nf=1.0 m=1
MP7 Y net6 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 net6 A6 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
.ends OA222X2_RVT




.subckt OA22X1_RVT A1 A2 A3 A4 VDD VSS Y
MP3 net3 A3 VDD VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP8 Y net6 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MN3 net6 A3 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net2 A1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 net6 A4 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends OA22X1_RVT




.subckt OA22X2_RVT A1 A2 A3 A4 VDD VSS Y
MP8 Y net6 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP4 net6 A4 net3 VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 net6 A4 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 Y net6 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 net6 A3 net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends OA22X2_RVT




.subckt OAI21X1_RVT A1 A2 A3 VDD VSS Y
MP3 net6 A3 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.46u l=0.03u nf=1.0 m=1
MP7 net7 net6 VDD VDD p105 w=0.17u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.46u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MN7 net7 net6 VSS VSS n105 w=0.10u l=0.03u nf=1.0 m=1
MN3 net6 A3 net2 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net2 A1 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
.ends OAI21X1_RVT




.subckt OAI21X2_RVT A1 A2 A3 VDD VSS Y
MP3 net6 A3 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP7 net7 net6 VDD VDD p105 w=0.26u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MN7 net7 net6 VSS VSS n105 w=0.16u l=0.03u nf=1.0 m=1
MN3 net6 A3 net2 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net2 A1 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.36u l=0.03u nf=1.0 m=1
.ends OAI21X2_RVT




.subckt OAI221X1_RVT A1 A2 A3 A4 A5 VDD VSS Y
MP5 net6 A5 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP7 net7 net6 VDD VDD p105 w=0.54u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net7 net6 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
.ends OAI221X1_RVT




.subckt OAI221X2_RVT A1 A2 A3 A4 A5 VDD VSS Y
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net7 net6 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP7 net7 net6 VDD VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP5 net6 A5 VDD VDD p105 w=0.19u l=0.03u nf=1.0 m=1
.ends OAI221X2_RVT




.subckt OAI222X1_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MP5 net5 A5 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 net6 A6 net5 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 net7 net6 VDD VDD p105 w=0.56u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 net6 A6 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 net7 net6 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
.ends OAI222X1_RVT




.subckt OAI222X2_RVT A1 A2 A3 A4 A5 A6 VDD VSS Y
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN7 net7 net6 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=1
MN3 net4 A3 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 net6 A6 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN4 net4 A4 net2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 net6 A5 net4 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP7 net7 net6 VDD VDD p105 w=0.75u l=0.03u nf=1.0 m=1
MP6 net6 A6 net5 VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP5 net5 A5 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
.ends OAI222X2_RVT




.subckt OAI22X1_RVT A1 A2 A3 A4 VDD VSS Y
MP3 net3 A3 VDD VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP7 net7 net6 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP8 Y net7 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MN7 net7 net6 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN3 net6 A3 net2 VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net2 A1 VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN4 net6 A4 net2 VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
.ends OAI22X1_RVT




.subckt OAI22X2_RVT A1 A2 A3 A4 VDD VSS Y
MP8 Y net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP7 net7 net6 VDD VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP4 net6 A4 net3 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP1 net1 A1 VDD VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP2 net6 A2 net1 VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MP3 net3 A3 VDD VDD p105 w=0.58u l=0.03u nf=1.0 m=1
MN2 net2 A2 VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN4 net6 A4 net2 VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN1 net2 A1 VSS VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN8 Y net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 net6 A3 net2 VSS n105 w=0.34u l=0.03u nf=1.0 m=1
MN7 net7 net6 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
.ends OAI22X2_RVT




.subckt OR2X1_RVT A1 A2 VDD VSS Y
MN0 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 SA1 A1 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MP0 Y SA1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP1 net95 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net95 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR2X1_RVT




.subckt OR2X2_RVT A1 A2 VDD VSS Y
MN0 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 SA1 A1 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MP0 Y SA1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net95 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net95 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR2X2_RVT




.subckt OR2X4_RVT A1 A2 VDD VSS Y
MN0 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN1 SA1 A1 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MP0 Y SA1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP1 net95 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 SA1 A2 net95 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR2X4_RVT




.subckt OR3X1_RVT A1 A2 A3 VDD VSS Y
MN1 SA1 A1 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN0 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN2 SA1 A2 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MP0 Y SA1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP1 net157 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net156 A2 net157 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 SA1 A3 net156 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR3X1_RVT




.subckt OR3X2_RVT A1 A2 A3 VDD VSS Y
MN1 SA1 A1 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN0 Y SA1 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN2 SA1 A2 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MP0 Y SA1 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net157 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net156 A2 net157 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 SA1 A3 net156 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR3X2_RVT




.subckt OR3X4_RVT A1 A2 A3 VDD VSS Y
MN4 SA2 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1 m=1
MN5 SA3 SA2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 SA1 A1 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN0 Y SA3 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN2 SA1 A2 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN3 SA1 A3 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MP4 SA2 SA1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP0 Y SA3 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP1 net176 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP2 net175 A2 net176 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP5 SA3 SA2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP3 SA1 A3 net175 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR3X4_RVT




.subckt OR4X1_RVT A1 A2 A3 A4 VDD VSS Y
MN5 net241 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1 m=1
MN6 net240 net241 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 SA1 A1 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN0 Y net240 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN3 SA1 A3 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN4 SA1 A4 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MP5 net241 SA1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP1 net239 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP0 Y net240 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP2 net238 A2 net239 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net237 A3 net238 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP6 net240 net241 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP4 SA1 A4 net237 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR4X1_RVT




.subckt OR4X2_RVT A1 A2 A3 A4 VDD VSS Y
MN5 net241 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1 m=1
MN6 net240 net241 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 SA1 A1 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN0 Y net240 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 SA1 A3 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN4 SA1 A4 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MP5 net241 SA1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP1 net239 A1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP0 Y net240 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP2 net238 A2 net239 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP3 net237 A3 net238 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP6 net240 net241 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP4 SA1 A4 net237 VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends OR4X2_RVT




.subckt OR4X4_RVT A1 A2 A3 A4 VDD VSS Y
MN5 net241 SA1 VSS VSS n105 w=0.21u l=0.03u nf=1 m=1
MN6 net240 net241 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 SA1 A1 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN2 SA1 A2 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN0 Y net240 VSS VSS n105 w=0.42u l=0.03u nf=1 m=4
MN3 SA1 A3 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MN4 SA1 A4 VSS VSS n105 w=0.13u l=0.03u nf=1.0 m=1
MP5 net241 SA1 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP1 net239 A1 VDD VDD p105 w=0.92u l=0.03u nf=1.0 m=1
MP0 Y net240 VDD VDD p105 w=0.8u l=0.03u nf=1 m=4
MP2 net238 A2 net239 VDD p105 w=0.92u l=0.03u nf=1.0 m=1
MP3 net237 A3 net238 VDD p105 w=0.92u l=0.03u nf=1.0 m=1
MP6 net240 net241 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP4 SA1 A4 net237 VDD p105 w=0.92u l=0.03u nf=1.0 m=1
.ends OR4X4_RVT



.GLOBAL VDD VSS
.subckt PGX1_RVT AN AP INOUT1 INOUT2 VDD VSS
MN INOUT1 AN INOUT2 VSS n105 w=0.375u l=0.03u nf=1 m=1
MP INOUT1 AP INOUT2 VDD p105 w=0.715u l=0.03u nf=1 m=1
.ends PGX1_RVT



.GLOBAL VDD VSS
.subckt PGX2_RVT AN AP INOUT1 INOUT2 VDD VSS
MN INOUT1 AN INOUT2 VSS n105 w=0.375u l=0.03u nf=1 m=2
MP INOUT1 AP INOUT2 VDD p105 w=0.715u l=0.03u nf=1 m=2
.ends PGX2_RVT



.GLOBAL VDD VSS
.subckt PGX4_RVT AN AP INOUT1 INOUT2 VDD VSS
MN INOUT1 AN INOUT2 VSS n105 w=0.375u l=0.03u nf=1 m=4
MP INOUT1 AP INOUT2 VDD p105 w=0.715u l=0.03u nf=1 m=4
.ends PGX4_RVT



.GLOBAL VDD
.subckt PMT1_RVT D G S VDD VSS
MP0 D G S VDD p105 w=0.8u l=0.03u nf=1 m=1
.ends PMT1_RVT



.GLOBAL VDD
.subckt PMT2_RVT D G S VDD VSS
MP0 D G S VDD p105 w=0.8u l=0.03u nf=1 m=2
.ends PMT2_RVT



.GLOBAL VDD
.subckt PMT3_RVT D G S VDD VSS
MP0 D G S VDD p105 w=0.8u l=0.03u nf=1 m=4
.ends PMT3_RVT




.subckt RDFFARX1_RVT CLK D Q QN RETN RSTB VDD VDDG VSS
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RDFFARX1_RVT




.subckt RDFFARX2_RVT CLK D Q QN RETN RSTB VDD VDDG VSS
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RDFFARX2_RVT




.subckt RDFFNARX1_RVT CLK D Q QN RETN RSTB VDD VDDG VSS
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RDFFNARX1_RVT




.subckt RDFFNARX2_RVT CLK D Q QN RETN RSTB VDD VDDG VSS
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RDFFNARX2_RVT




.subckt RDFFNSRARX1_RVT CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRARX1_RVT




.subckt RDFFNSRARX2_RVT CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRARX2_RVT




.subckt RDFFNSRASRNX1_RVT CLK D NRESTORE QN RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASRNX1_RVT




.subckt RDFFNSRASRNX2_RVT CLK D NRESTORE QN RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASRNX2_RVT




.subckt RDFFNSRASRQX1_RVT CLK D NRESTORE Q RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASRQX1_RVT




.subckt RDFFNSRASRQX2_RVT CLK D NRESTORE Q RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASRQX2_RVT




.subckt RDFFNSRASRX1_RVT CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASRX1_RVT




.subckt RDFFNSRASRX2_RVT CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASRX2_RVT




.subckt RDFFNSRASX1_RVT CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM2 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASX1_RVT




.subckt RDFFNSRASX2_RVT CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM2 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFNSRASX2_RVT




.subckt RDFFNSRX1_RVT CLK D NRESTORE Q QN SAVE VDD VDDG VSS
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn1 net403 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net400 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net366 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net366 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM11 net403 net400 net390 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM3 net400 net403 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM12 net390 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM14 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net400 net403 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net400 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net403 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM4 net363 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net363 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM9 net403 net400 net391 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM10 net391 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends RDFFNSRX1_RVT




.subckt RDFFNSRX2_RVT CLK D NRESTORE Q QN SAVE VDD VDDG VSS
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn1 net403 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net400 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net366 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net366 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM11 net403 net400 net390 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM3 net400 net403 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM12 net390 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM14 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net400 net403 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net400 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net403 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM4 net363 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net363 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM9 net403 net400 net391 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM10 net391 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends RDFFNSRX2_RVT




.subckt RDFFNX1_RVT CLK D Q QN RETN VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
.ends RDFFNX1_RVT




.subckt RDFFNX2_RVT CLK D Q QN RETN VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
.ends RDFFNX2_RVT




.subckt RDFFSRARX1_RVT CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRARX1_RVT




.subckt RDFFSRARX2_RVT CLK D NRESTORE Q QN RSTB SAVE VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRARX2_RVT




.subckt RDFFSRASRX1_RVT CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRASRX1_RVT




.subckt RDFFSRASRX2_RVT CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRASRX2_RVT




.subckt RDFFSRASX1_RVT CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM2 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRASX1_RVT




.subckt RDFFSRASX2_RVT CLK D NRESTORE Q QN SAVE SETB VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM2 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRASX2_RVT




.subckt RDFFSRSSRX1_RVT CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn16 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn23 rrr SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 rrr D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 Q net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 QN net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp17 rrr RSTB net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 net01 SET VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp16 rrr D net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 VDD net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 QN net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 Q net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRSSRX1_RVT




.subckt RDFFSRSSRX2_RVT CLK D NRESTORE Q QN RSTB SAVE SETB VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn16 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn23 rrr SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 rrr D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 Q net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 QN net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp17 rrr RSTB net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 net01 SET VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp16 rrr D net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 VDD net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 QN net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 Q net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RDFFSRSSRX2_RVT




.subckt RDFFSRX1_RVT CLK D NRESTORE Q QN SAVE VDD VDDG VSS
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn1 net403 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net400 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net366 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net366 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM11 net403 net400 net390 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM3 net400 net403 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM12 net390 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM14 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net400 net403 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net400 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net403 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM4 net363 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net363 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM9 net403 net400 net391 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM10 net391 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends RDFFSRX1_RVT




.subckt RDFFSRX2_RVT CLK D NRESTORE Q QN SAVE VDD VDDG VSS
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn1 net403 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net400 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net366 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net366 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf D VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM11 net403 net400 net390 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM3 net400 net403 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM12 net390 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM14 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net400 net403 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net400 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net403 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM4 net363 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net363 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf D VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM9 net403 net400 net391 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM10 net391 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
.ends RDFFSRX2_RVT




.subckt RDFFX1_RVT CLK D Q QN RETN VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP2 netp2 D netp1 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
.ends RDFFX1_RVT




.subckt RDFFX2_RVT CLK D Q QN RETN VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 D netn1 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP2 netp2 D netp1 VDD p105 w=0.45u l=0.03u nf=1 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.45u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
.ends RDFFX2_RVT




.subckt RSDFFARX1_RVT CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
MN01 INP INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 INP netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP01 INP INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 INP netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RSDFFARX1_RVT




.subckt RSDFFARX2_RVT CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
MN01 INP INN VSS VSS n105 w=0.389u l=0.03u nf=1.0 m=1
MN05 INN SI netn04 VSS n105 w=0.389u l=0.03u nf=1.0 m=1
MN04 netn04 SE VSS VSS n105 w=0.389u l=0.03u nf=1.0 m=1
MN02 netn02 SEN VSS VSS n105 w=0.389u l=0.03u nf=1.0 m=1
MN03 INN D netn02 VSS n105 w=0.389u l=0.03u nf=1.0 m=1
MNSE SEN SE VSS VSS n105 w=0.389u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 INP netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP01 INP INN VDD VDD p105 w=0.724u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.724u l=0.03u nf=1.0 m=1
MP05 INN SI netp04 VDD p105 w=0.724u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.724u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.724u l=0.03u nf=1.0 m=1
MPSE SEN SE VDD VDD p105 w=0.724u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 INP netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RSDFFARX2_RVT




.subckt RSDFFNARX1_RVT CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
MN01 INP INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 INP netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP01 INP INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 INP netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RSDFFNARX1_RVT




.subckt RSDFFNARX2_RVT CLK D Q QN RETN RSTB SE SI VDD VDDG VSS
MN01 INP INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNR1 r RSTB VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN15 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 net336 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 net336 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN4 netp4 r VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN2 netp2 INP netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP01 INP INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPR1 r RSTB VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP15 netp26 netp22 netp25 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP14 netp25 r VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP3 netp3 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 netp4 r netp3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP2 netp2 INP netp1 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1.0 m=1
.ends RSDFFNARX2_RVT




.subckt RSDFFNSRARX1_RVT CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRARX1_RVT




.subckt RSDFFNSRARX2_RVT CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRARX2_RVT




.subckt RSDFFNSRASRNX1_RVT CLK D NRESTORE QN RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASRNX1_RVT




.subckt RSDFFNSRASRNX2_RVT CLK D NRESTORE QN RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASRNX2_RVT




.subckt RSDFFNSRASRQX1_RVT CLK D NRESTORE Q RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASRQX1_RVT




.subckt RSDFFNSRASRQX2_RVT CLK D NRESTORE Q RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASRQX2_RVT




.subckt RSDFFNSRASRX1_RVT CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASRX1_RVT




.subckt RSDFFNSRASRX2_RVT CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASRX2_RVT




.subckt RSDFFNSRASX1_RVT CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM47 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM45 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM43 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM42 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM41 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM40 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM49 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM44 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM39 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM38 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM2 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASX1_RVT




.subckt RSDFFNSRASX2_RVT CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM47 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM45 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM43 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM42 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM41 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM40 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKP hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM49 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM44 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM39 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM38 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM2 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRASX2_RVT




.subckt RSDFFNSRX1_RVT CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
MM8 net1556 net8 net346 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net346 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net356 CLKP hjf VSS n105 w=0.35u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net356 net2 net342 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM1 net2 net356 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM3 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn4 net342 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net356 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net2 net356 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp6 net356 net2 net360 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net360 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRX1_RVT




.subckt RSDFFNSRX2_RVT CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
MM8 net1556 net8 net346 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net346 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKN _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net356 CLKP hjf VSS n105 w=0.35u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net356 net2 net342 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM1 net2 net356 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM3 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn4 net342 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKP _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net356 CLKN hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net2 net356 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp6 net356 net2 net360 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net360 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFNSRX2_RVT




.subckt RSDFFNX1_RVT CLK D Q QN RETN SE SI VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 net373 netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN01 net373 INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP2 netp2 net373 netp1 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 net373 INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
.ends RSDFFNX1_RVT




.subckt RSDFFNX2_RVT CLK D Q QN RETN SE SI VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKP netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 net336 netn1 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN1 netn1 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN01 net336 INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP5 netp5 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP12 netp8 CLKN netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKP VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP2 netp2 net336 netp1 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP1 netp1 CLKN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 net336 INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
.ends RSDFFNX2_RVT




.subckt RSDFFSRARX1_RVT CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRARX1_RVT




.subckt RSDFFSRARX2_RVT CLK D NRESTORE Q QN RSTB SAVE SE SI VDD VDDG VSS
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRARX2_RVT




.subckt RSDFFSRASRX1_RVT CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRASRX1_RVT




.subckt RSDFFSRASRX2_RVT CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
Mmn29 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn12 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn10 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn28 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn27 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 RSTB _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmp29 net1556 SETB net444 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
Mmp12 net1556 net8 net444 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
Mmp10 net444 CLKP VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
Mmp28 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp27 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRASRX2_RVT




.subckt RSDFFSRASX1_RVT CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM47 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM45 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM43 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM42 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM41 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM40 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM49 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM44 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM39 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM38 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM2 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRASX1_RVT




.subckt RSDFFSRASX2_RVT CLK D NRESTORE Q QN SAVE SE SETB SI VDD VDDG VSS
MM66 net1556 net8 _n1247 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM64 _n1247 SETB _n1248 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM63 _n1248 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM60 net994 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM58 net2 SETB net994 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM47 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM45 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM43 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM42 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM41 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM40 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM37 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM33 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM32 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM30 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM23 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM22 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM21 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM19 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM16 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM15 net155 net2 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM11 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM9 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM8 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM3 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM57 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM56 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM51 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM50 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM36 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM28 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
MM55 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM54 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM53 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM52 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM35 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM27 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM67 net1556 SETB net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM65 net1556 net8 net444 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM62 net444 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM61 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM59 net2 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM49 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM44 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM39 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM38 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM34 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM31 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM29 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM26 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM25 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM24 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM20 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM18 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM17 net155 VDD net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM14 net155 net2 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM12 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM10 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM7 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM5 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM2 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRASX2_RVT




.subckt RSDFFSRSSRX1_RVT CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
MN05 net04 SI VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN01 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN02 net02 SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN07 net05 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN06 hjf net05 net02 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN08 hjf SE net04 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN03 net02 D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn5 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MP05 net04 SI VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP04 net02 RSTB net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP07 net05 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP08 hjf net05 net04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP06 hjf SE net02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP01 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 net02 D net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 net01 SET VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 VDD net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends RSDFFSRSSRX1_RVT




.subckt RSDFFSRSSRX2_RVT CLK D NRESTORE Q QN RSTB SAVE SE SETB SI VDD VDDG VSS
MN05 net04 SI VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN01 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM3 net358 net155 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net341 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN02 net02 SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM5 net341 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN07 net05 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN06 hjf net05 net02 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN08 hjf SE net04 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN03 net02 D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net358 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net155 CLKN hjf VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net155 net358 _n989 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn8 net9 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn9 net8 VDD net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn5 _n989 VDD _n991 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn4 _n991 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MP05 net04 SI VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM2 net358 net155 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP04 net02 RSTB net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP07 net05 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP08 hjf net05 net04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM6 net1556 net8 net347 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP06 hjf SE net02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM4 net347 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP01 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 net02 D net01 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 net01 SET VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net358 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net155 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp9 net8 VDD VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp5 net155 VDD net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp6 net155 net358 net348 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp8 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net348 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
.ends RSDFFSRSSRX2_RVT




.subckt RSDFFSRX1_RVT CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
MM8 net1556 net8 net346 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net346 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net356 CLKN hjf VSS n105 w=0.35u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn6 net356 net2 net342 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM1 net2 net356 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM3 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
Mmn4 net342 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net356 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net2 net356 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp6 net356 net2 net360 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net360 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRX1_RVT




.subckt RSDFFSRX2_RVT CLK D NRESTORE Q QN SAVE SE SI VDD VDDG VSS
MM8 net1556 net8 net346 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM6 net346 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn25 p1 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn24 rrr _n53 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn23 _n53 D _n52 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn17 _n53 SI net6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn16 net6 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn3 _n52 p1 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmn26 RESTORE NRESTORE VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn18 _n766 jk netn10 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn19 netn10 RESTORE VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM0 net2 NRESTORE _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn7 net1556 CLKP _n766 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn1 net356 CLKN hjf VSS n105 w=0.35u l=0.03u nf=1.0 m=1
Mmn012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn14 QN net1556 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn6 net356 net2 net342 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM1 net2 net356 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MM3 net8 net1556 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
Mmn13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
Mmn4 net342 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
Mmn03 hjf rrr VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
Mmp32 netp103 SAVEN VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp33 jk2 net8 netp103 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp21 jk2 jk netp102 VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp20 netp102 SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp22 SAVEN SAVE VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmp15 jk jk2 VDDG VDDG p105_hvt w=0.4u l=0.03u nf=1.0 m=1
Mmn33 jk2 net8 netn103 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn32 netn103 SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn20 jk2 jk netn102 VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn21 netn102 SAVEN VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn22 SAVEN SAVE VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
Mmn15 jk jk2 VSS VSS n105_hvt w=0.3u l=0.03u nf=1.0 m=1
MM7 net1556 net8 net4 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM5 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp25 _n53 SI net5 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp24 p1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp23 rrr _n53 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp17 net5 p1 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp16 _n53 D _n50 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp3 _n50 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
Mmp26 RESTORE NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp18 netp10 NRESTORE VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp19 _n766 jk netp10 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp11 net2 RESTORE _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp7 net1556 CLKN _n766 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp1 net356 CLKP hjf VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MM2 net2 net356 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp6 net356 net2 net360 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM4 net8 net1556 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
Mmp13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
Mmp4 net360 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
Mmp14 QN net1556 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
Mmp03 hjf rrr VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFSRX2_RVT




.subckt RSDFFX1_RVT CLK D Q QN RETN SE SI VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 INP netn1 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN01 INP INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=1
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.4u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP2 netp2 INP netp1 VDD p105 w=0.45u l=0.03u nf=1 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.45u l=0.03u nf=1 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 INP INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFX1_RVT




.subckt RSDFFX2_RVT CLK D Q QN RETN SE SI VDD VDDG VSS
MN3 netp4 netp2 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN14 netp26 netp22 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN6 netp2 netp4 netn5 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN5 netn5 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN12 netp8 CLKN netp27 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN13 netp27 netp26 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN20 netp20 RETN VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN16 netn23 RETN VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN19 netp22 DL netn23 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN18 netn21 netp20 VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN17 netp22 QL netn21 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN10 Q netp8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN11 QN DL VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN9 DL netp8 VSS VSS n105 w=0.40u l=0.03u nf=1 m=1
MN7 netn7 CLKP VSS VSS n105 w=0.30u l=0.03u nf=1 m=1
MN8 netp8 netp4 netn7 VSS n105 w=0.30u l=0.03u nf=1 m=1
MN2 netp2 INP netn1 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN1 netn1 CLKN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN02 netn02 SEN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN05 INN SI netn04 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN04 netn04 SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN01 INP INN VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MNSE SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1 m=1
MN03 INN D netn02 VSS n105 w=0.25u l=0.03u nf=1 m=1
MN21 RETNN RETN VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN25 netp102 RETNN QL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN24 QL netp103 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN23 netp103 netp102 VSS VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MN22 netp102 RETN DL VSS n105_hvt w=0.30u l=0.03u nf=1 m=1
MP25 netp102 RETN QL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP24 QL netp103 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP23 netp103 netp102 VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP21 RETNN RETN VDDG VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP22 netp102 RETNN DL VDDG p105_hvt w=0.40u l=0.03u nf=1 m=1
MP3 netp4 netp2 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1 m=1
MP6 netp2 netp4 netp5 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP5 netp5 CLKN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP12 netp8 CLKP netp27 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP13 netp27 netp26 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP14 netp26 netp22 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP20 netp20 RETN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP18 netp23 netp20 VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP19 netp22 DL netp23 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP17 netp22 QL netp21 VDD p105 w=0.30u l=0.03u nf=1 m=1
MP16 netp21 RETN VDD VDD p105 w=0.30u l=0.03u nf=1 m=1
MP10 Q netp8 VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP11 QN DL VDD VDD p105 w=0.80u l=0.03u nf=1 m=2
MP9 DL netp8 VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP7 netp7 CLKN VDD VDD p105 w=0.40u l=0.03u nf=1 m=1
MP8 netp8 netp4 netp7 VDD p105 w=0.40u l=0.03u nf=1 m=1
MP2 netp2 INP netp1 VDD p105 w=0.45u l=0.03u nf=1 m=1
MP1 netp1 CLKP VDD VDD p105 w=0.45u l=0.03u nf=1 m=1
MP05 INN SI netp04 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 netp04 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 INP INN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MPSE SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 INN D netp02 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 netp02 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends RSDFFX2_RVT




.subckt SDFFARX1_RVT CLK D Q QN RSTB SE SI VDD VSS
MN8 net293 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN02 SA2 SEN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net293 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
.ends SDFFARX1_RVT




.subckt SDFFARX2_RVT CLK D Q QN RSTB SE SI VDD VSS
MN8 net293 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN02 SA2 SEN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net293 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
.ends SDFFARX2_RVT



.GLOBAL VDD
.subckt SDFFASRSX1_RVT CLK D Q QN RSTB SE SETB SI SO VDD VSS
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP6 D2 D3 FB1 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP15 SO D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net388 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 D3 SETB net390 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 net388 D4 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN6 D2 D3 FB2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net390 D2 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN15 SO D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFASRSX1_RVT




.subckt SDFFASRSX2_RVT CLK D Q QN RSTB SE SETB SI SO VDD VSS
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP6 D2 D3 FB1 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP15 SO D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net388 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 D3 SETB net389 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 net388 D4 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN6 D2 D3 FB2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN2 net389 D2 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.2u l=0.03u nf=1.0 m=1
MN1 D1 CLKN D2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN15 SO D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFASRSX2_RVT




.subckt SDFFASRX1_RVT CLK D Q QN RSTB SE SETB SI VDD VSS
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP13 Q D5 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 D3 SETB net253 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net252 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN8 net252 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net253 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends SDFFASRX1_RVT




.subckt SDFFASRX2_RVT CLK D Q QN RSTB SE SETB SI VDD VSS
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD D4 D5 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 D5 RSTB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 RSTB FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN3 D3 SETB net253 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 D5 RSTB net252 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN4 FB3 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 FB2 RSTB FB3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN8 net252 D4 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net253 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends SDFFASRX2_RVT




.subckt SDFFASX1_RVT CLK D Q QN SE SETB SI VDD VSS
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 D5 D4 VSS VSS n105 w=0.27u l=0.03u nf=1 m=1
MN3 D3 SETB net242 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net242 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP8 D5 D4 VDD VDD p105 w=0.76u l=0.03u nf=1.0 m=1
.ends SDFFASX1_RVT




.subckt SDFFASX2_RVT CLK D Q QN SE SETB SI VDD VSS
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 D5 D4 VSS VSS n105 w=0.27u l=0.03u nf=1 m=1
MN3 D3 SETB net242 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN12 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 FB6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 FB5 SETB FB6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 net242 D2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 SETB FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP3 D3 SETB VDD VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MP12 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP2 VDD D2 D3 VDD p105 w=0.52u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP8 D5 D4 VDD VDD p105 w=0.76u l=0.03u nf=1.0 m=1
.ends SDFFASX2_RVT




.subckt SDFFNARX1_RVT CLK D Q QN RSTB SE SI VDD VSS
MM19 VDD net7 net227 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net227 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP26 VDD net228 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net228 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net2 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net7 CLKN net230 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net228 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 net228 CLKP net227 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM45 net234 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 net229 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 net230 D net229 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM52 net230 SI net232 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM53 net232 net234 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM18 net227 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net227 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM49 net231 net234 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM50 net233 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN25 net3 net228 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN23 net228 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net228 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net7 CLKP net230 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN7 net228 CLKN net227 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM47 net230 D net231 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM44 net234 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM51 net230 SI net233 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFNARX1_RVT




.subckt SDFFNARX2_RVT CLK D Q QN RSTB SE SI VDD VSS
MM19 VDD net7 net227 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP16 net7 net227 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP15 net7 RSTB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP8 net10 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP27 net2 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP26 VDD net228 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net228 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net2 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net7 CLKN net230 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP21 net4 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP20 net228 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP7 net228 CLKP net227 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM45 net234 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 net229 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 net230 D net229 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM52 net230 SI net232 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM53 net232 net234 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM18 net227 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN17 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 net11 RSTB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 net7 net227 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM49 net231 net234 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM50 net233 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN25 net3 net228 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN23 net228 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN net228 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net2 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net7 CLKP net230 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN22 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN24 net2 RSTB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN7 net228 CLKN net227 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM47 net230 D net231 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM44 net234 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM51 net230 SI net233 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFNARX2_RVT




.subckt SDFFNASRX1_RVT CLK D Q QN RSTB SE SETB SI VDD VSS
MM51 net01 SI net211 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM44 net212 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM47 net01 D net209 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM49 net209 net212 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM50 net211 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM52 net01 SI net210 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM53 net210 net212 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM45 net212 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 net01 D net208 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 net208 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends SDFFNASRX1_RVT




.subckt SDFFNASRX2_RVT CLK D Q QN RSTB SE SETB SI VDD VSS
MM51 net01 SI net211 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM44 net212 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM47 net01 D net209 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM49 net209 net212 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM50 net211 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN5 net5 RSTB net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 net1 net2 net5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net9 net7 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN9 net8 RSTB net9 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM52 net01 SI net210 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM53 net210 net212 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM45 net212 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM46 net01 D net208 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 net208 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP5 net1 RSTB net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP9 net8 RSTB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 net8 net7 VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP4 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
.ends SDFFNASRX2_RVT




.subckt SDFFNASX1_RVT CLK D Q QN SE SETB SI VDD VSS
MM12 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM11 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD net7 net8 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP16 net01 D net184 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP22 net01 SI net186 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP15 net188 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP18 net184 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP23 net186 net188 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM14 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net8 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN21 net01 SI net187 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN20 net187 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN19 net185 net188 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN15 net188 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN17 net01 D net185 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFNASX1_RVT




.subckt SDFFNASX2_RVT CLK D Q QN SE SETB SI VDD VSS
MM12 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM11 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP3 net2 SETB VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 VDD net1 net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP8 VDD net7 net8 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MP14 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net1 CLKN net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP12 net7 net8 net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP11 net7 SETB net10 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP10 net10 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP16 net01 D net184 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP22 net01 SI net186 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP15 net188 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP18 net184 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP23 net186 net188 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM14 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM13 net6 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net3 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN3 net2 SETB net3 VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN8 net8 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN14 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 net1 CLKP net01 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN10 net12 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 net11 SETB net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 net7 net8 net11 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN21 net01 SI net187 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN20 net187 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN19 net185 net188 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN15 net188 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN17 net01 D net185 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFNASX2_RVT




.subckt SDFFNX1_RVT CLK D Q QN SE SI VDD VSS
MM28 net7 net268 net269 VDD p105 w=0.3u l=0.03u nf=1 m=1
MM27 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM25 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM24 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MM39 VDD net7 net268 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MM37 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM35 Q net268 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MM32 net1 CLKN net277 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM41 VDD net1 net2 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MM29 net269 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM52 net277 SI net274 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM53 net274 net276 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM45 net276 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM55 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM57 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM46 net277 D net272 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 net272 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM26 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM38 net268 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MM36 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MM34 Q net268 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MM33 net1 CLKP net277 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM31 net270 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM42 net1 net2 net271 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM30 net271 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM40 net2 net1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MM51 net277 SI net275 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM43 net7 net268 net270 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM44 net276 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM54 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM56 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM47 net277 D net273 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM49 net273 net276 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM50 net275 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFNX1_RVT




.subckt SDFFNX2_RVT CLK D Q QN SE SI VDD VSS
MM28 net7 net268 net269 VDD p105 w=0.3u l=0.03u nf=1 m=1
MM27 net7 CLKP net2 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM25 net4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM24 net1 net2 net4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MM39 VDD net7 net268 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MM37 QN net7 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM35 Q net268 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MM32 net1 CLKN net277 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MM41 VDD net1 net2 VDD p105 w=0.7u l=0.03u nf=1.0 m=1
MM29 net269 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MM52 net277 SI net274 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM53 net274 net276 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM45 net276 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM55 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM57 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MM46 net277 D net272 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM48 net272 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MM26 net7 CLKN net2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM38 net268 net7 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MM36 QN net7 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM34 Q net268 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MM33 net1 CLKP net277 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM31 net270 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM42 net1 net2 net271 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM30 net271 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM40 net2 net1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MM51 net277 SI net275 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM43 net7 net268 net270 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MM44 net276 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM54 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM56 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MM47 net277 D net273 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM49 net273 net276 VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MM50 net275 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFNX2_RVT



.GLOBAL VDD VSS
.subckt SDFFSSRX1_RVT CLK D Q QN RSTB SE SETB SI VDD VSS
MN6 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN05 net04 SI VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN01 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN08 net06 SE net04 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN07 net05 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN06 net06 net05 net02 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 net02 SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN03 net02 D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 IQN net8 net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 net1 CLKN net06 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 IQN CLKP net2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN IQN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN8 net8 IQN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net2 net1 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP05 net04 SI VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP08 net06 net05 net04 VDD p105 w=0.35u l=0.03u nf=1.0 m=1
MP07 net05 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP06 net06 SE net02 VDD p105 w=0.35u l=0.03u nf=1.0 m=1
MP04 net02 RSTB net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP03 net02 D net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP02 net01 SET VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP10 net10 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP12 IQN net8 net10 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 net1 CLKP net06 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 IQN CLKN net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP4 net4 CLKN VDD VDD p105 w=0.25u l=0.03u nf=1.0 m=1
MP14 QN IQN VDD VDD p105 w=0.8u l=0.03u nf=1 m=1
MP8 net8 IQN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFSSRX1_RVT




.subckt SDFFSSRX2_RVT CLK D Q QN RSTB SE SETB SI VDD VSS
MN6 net1 net2 net6 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 net2 net1 VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN13 Q net8 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN05 net04 SI VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN01 SET SETB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN08 net06 SE net04 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN07 net05 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN06 net06 net05 net02 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 net02 SET net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN03 net02 D net03 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 net03 RSTB VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 net12 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN12 IQN net8 net12 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 net6 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 net1 CLKN net06 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 IQN CLKP net2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN14 QN IQN VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN8 net8 IQN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN012 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MN011 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net2 net1 VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP13 Q net8 VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP05 net04 SI VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP01 SET SETB VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP08 net06 net05 net04 VDD p105 w=0.35u l=0.03u nf=1.0 m=1
MP07 net05 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP06 net06 SE net02 VDD p105 w=0.35u l=0.03u nf=1.0 m=1
MP04 net02 RSTB net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP03 net02 D net01 VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP02 net01 SET VDD VDD p105 w=0.6u l=0.03u nf=1.0 m=1
MP10 net10 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP12 IQN net8 net10 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP1 net1 CLKP net06 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP7 IQN CLKN net2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP4 net4 CLKN VDD VDD p105 w=0.25u l=0.03u nf=1.0 m=1
MP14 QN IQN VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP8 net8 IQN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP012 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP011 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP6 net1 net2 net4 VDD p105 w=0.25u l=0.03u nf=1.0 m=1
.ends SDFFSSRX2_RVT




.subckt SDFFX1_RVT CLK D Q QN SE SI VDD VSS
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP12 D5 D4 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 D5 D4 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=1
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends SDFFX1_RVT




.subckt SDFFX2_RVT CLK D Q QN SE SI VDD VSS
MP4 FB1 CLKN VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MPC1 CLKN CLK VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MPC2 CLKP CLKN VDD VDD p105 w=0.74u l=0.03u nf=1.0 m=1
MP1 D1 CLKP D2 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP01 SEN SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP10 FB4 CLKP VDD VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 D3 D2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP03 D1 D SA1 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP02 SA1 SE VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP05 D1 SI SA3 VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP04 SA3 SEN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP12 D5 D4 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP14 QN D4 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP13 Q D5 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP7 D4 CLKN D3 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP11 D4 D5 FB4 VDD p105 w=0.3u l=0.03u nf=1 m=1
MP5 D2 D3 FB1 VDD p105 w=0.3u l=0.03u nf=1 m=1
MNC1 CLKN CLK VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MNC2 CLKP CLKN VSS VSS n105 w=0.4u l=0.03u nf=1 m=1
MN2 D3 D2 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN01 SEN SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN12 D5 D4 VSS VSS n105 w=0.35u l=0.03u nf=1 m=1
MN10 FB5 CLKN VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN03 D1 D SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN02 SA2 SEN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN04 SA4 SE VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN05 D1 SI SA4 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN14 QN D4 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN13 Q D5 VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN1 D1 CLKN D2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN7 D4 CLKP D3 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 D2 D3 FB2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN4 FB2 CLKP VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN11 D4 D5 FB5 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
.ends SDFFX2_RVT




.subckt SHFILL128_RVT VDD VSS
.ends SHFILL128_RVT




.subckt SHFILL1_RVT VDD VSS
.ends SHFILL1_RVT




.subckt SHFILL2_RVT VDD VSS
.ends SHFILL2_RVT




.subckt SHFILL3_RVT VDD VSS
.ends SHFILL3_RVT




.subckt SHFILL64_RVT VDD VSS
.ends SHFILL64_RVT




.subckt TIEH_RVT VDD VSS Y
MN0 net47 net47 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP0 Y net47 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends TIEH_RVT




.subckt TIEL_RVT VDD VSS Y
MN0 Y net42 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP0 net42 net42 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends TIEL_RVT




.subckt TNBUFFX16_RVT A EN VDD VSS Y
MN5 Y net128 VSS VSS n105 w=0.375u l=0.03u nf=1 m=16
MN4 VSS net126 net128 VSS n105 w=0.38u l=0.03u nf=1 m=3
MN2 net128 A VSS VSS n105 w=0.42u l=0.03u nf=1 m=3
MN3 net127 EN net128 VSS n105 w=0.43u l=0.03u nf=1 m=3
MN1 net126 EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MP5 Y net127 VDD VDD p105 w=0.715u l=0.03u nf=1 m=16
MP4 net127 net126 net128 VDD p105 w=0.55u l=0.03u nf=1 m=3
MP3 VDD EN net127 VDD p105 w=0.55u l=0.03u nf=1 m=3
MP2 net127 A VDD VDD p105 w=0.8u l=0.03u nf=1 m=3
MP1 net126 EN VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
.ends TNBUFFX16_RVT




.subckt TNBUFFX1_RVT A EN VDD VSS Y
MN5 Y net128 VSS VSS n105 w=0.375u l=0.03u nf=1.0 m=1
MN4 VSS net126 net128 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 net128 A VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 net127 EN net128 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN1 net126 EN VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MP5 Y net127 VDD VDD p105 w=0.715u l=0.03u nf=1.0 m=1
MP4 net127 net126 net128 VDD p105 w=0.25u l=0.03u nf=1.0 m=1
MP3 VDD EN net127 VDD p105 w=0.3u l=0.03u nf=1.0 m=1
MP2 net127 A VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP1 net126 EN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
.ends TNBUFFX1_RVT




.subckt TNBUFFX2_RVT A EN VDD VSS Y
MN5 Y net128 VSS VSS n105 w=0.375u l=0.03u nf=1 m=2
MN4 VSS net126 net128 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN2 net128 A VSS VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN3 net127 EN net128 VSS n105 w=0.26u l=0.03u nf=1.0 m=1
MN1 net126 EN VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MP5 Y net127 VDD VDD p105 w=0.715u l=0.03u nf=1 m=2
MP4 net127 net126 net128 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP3 VDD EN net127 VDD p105 w=0.4u l=0.03u nf=1.0 m=1
MP2 net127 A VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP1 net126 EN VDD VDD p105 w=0.4u l=0.03u nf=1.0 m=1
.ends TNBUFFX2_RVT




.subckt TNBUFFX32_RVT A EN VDD VSS Y
MN6 net175 A VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN0 net173 EN VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN7 net174 net175 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN5 Y net171 VSS VSS n105 w=0.375u l=0.03u nf=1 m=32
MN4 VSS net173 net171 VSS n105 w=0.38u l=0.03u nf=1 m=6
MN2 net171 net174 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=6
MN3 net170 net172 net171 VSS n105 w=0.43u l=0.03u nf=1.0 m=6
MN1 net172 net173 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MP6 net175 A VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
MP7 net174 net175 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP0 net173 EN VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP5 Y net170 VDD VDD p105 w=0.715u l=0.03u nf=1 m=32
MP4 net170 net173 net171 VDD p105 w=0.55u l=0.03u nf=1 m=6
MP3 VDD net172 net170 VDD p105 w=0.55u l=0.03u nf=1 m=6
MP2 net170 net174 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=6
MP1 net172 net173 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
.ends TNBUFFX32_RVT




.subckt TNBUFFX4_RVT A EN VDD VSS Y
MN5 Y net128 VSS VSS n105 w=0.375u l=0.03u nf=1 m=4
MN4 VSS net126 net128 VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN2 net128 A VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN3 net127 EN net128 VSS n105 w=0.43u l=0.03u nf=1.0 m=1
MN1 net126 EN VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MP5 Y net127 VDD VDD p105 w=0.715u l=0.03u nf=1 m=4
MP4 net127 net126 net128 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP3 VDD EN net127 VDD p105 w=0.55u l=0.03u nf=1.0 m=1
MP2 net127 A VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP1 net126 EN VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
.ends TNBUFFX4_RVT




.subckt TNBUFFX8_RVT A EN VDD VSS Y
MN5 Y net128 VSS VSS n105 w=0.375u l=0.03u nf=1 m=8
MN4 VSS net126 net128 VSS n105 w=0.38u l=0.03u nf=1 m=2
MN2 net128 A VSS VSS n105 w=0.42u l=0.03u nf=1 m=2
MN3 net127 EN net128 VSS n105 w=0.43u l=0.03u nf=1 m=2
MN1 net126 EN VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MP5 Y net127 VDD VDD p105 w=0.715u l=0.03u nf=1 m=8
MP4 net127 net126 net128 VDD p105 w=0.55u l=0.03u nf=1 m=2
MP3 VDD EN net127 VDD p105 w=0.55u l=0.03u nf=1 m=2
MP2 net127 A VDD VDD p105 w=0.8u l=0.03u nf=1 m=2
MP1 net126 EN VDD VDD p105 w=0.5u l=0.03u nf=1.0 m=1
.ends TNBUFFX8_RVT




.subckt XNOR2X1_RVT A1 A2 VDD VSS Y
MN2 A2B A2 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN5 Y1 A1 SA4 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN1 A1B A1 VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN7 Y Y1 VSS VSS n105 w=0.41u l=0.03u nf=1.0 m=1
MN4 SA2 A2B VSS VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MN3 Y1 A1B SA2 VSS n105 w=0.22u l=0.03u nf=1.0 m=1
MP2 A2B A2 VDD VDD p105 w=0.44u l=0.03u nf=1.0 m=1
MP7 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 A1B A1 VDD VDD p105 w=0.44u l=0.03u nf=1.0 m=1
MP6 Y1 A1 SA3 VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.47u l=0.03u nf=1.0 m=1
MP4 Y1 A1B SA1 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
.ends XNOR2X1_RVT




.subckt XNOR2X2_RVT A1 A2 VDD VSS Y
MN7 Y Y1 VSS VSS n105 w=0.40u l=0.03u nf=1.0 m=2
MN1 A1B A1 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN5 Y1 A1 SA4 VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN3 Y1 A1B SA2 VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN4 SA2 A2B VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP2 A2B A2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP6 Y1 A1 SA3 VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP1 A1B A1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP7 Y Y1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP4 Y1 A1B SA1 VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
.ends XNOR2X2_RVT




.subckt XNOR3X1_RVT A1 A2 A3 VDD VSS Y
MN4 SA2 A2B VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN8 Y1B Y1 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 A1B A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.40u l=0.03u nf=1.0 m=1
MN5 Y1 A1 SA4 VSS n105 w=0.40u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 A3B A3 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN11 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN9 Y1 A3B Y2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN3 Y1 A1B SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=1
MN10 Y1B A3 Y2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MP2 A2B A2 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP6 Y1 A1 SA3 VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP11 Y Y2 VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=1
MP8 Y1B Y1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP7 A3B A3 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP4 Y1 A1B SA1 VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP10 Y1B A3B Y2 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.65u l=0.03u nf=1.0 m=1
MP1 A1B A1 VDD VDD p105 w=0.50u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP9 Y1 A3 Y2 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
.ends XNOR3X1_RVT




.subckt XNOR3X2_RVT A1 A2 A3 VDD VSS Y
MP10 Y1B A3B Y2 VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP4 Y1 A1B SA1 VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP7 A3B A3 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP8 Y1B Y1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP11 Y Y2 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=2
MP2 A2B A2 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP6 Y1 A1 SA3 VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP9 Y1 A3 Y2 VDD p105 w=0.38u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MP1 A1B A1 VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=1
MN11 Y Y2 VSS VSS n105 w=0.40u l=0.03u nf=1.0 m=2
MN1 A1B A1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN7 A3B A3 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN8 Y1B Y1 VSS VSS n105 w=0.30u l=0.03u nf=1.0 m=1
MN4 SA2 A2B VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN5 Y1 A1 SA4 VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN10 Y1B A3 Y2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN3 Y1 A1B SA2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN9 Y1 A3B Y2 VSS n105 w=0.35u l=0.03u nf=1.0 m=1
.ends XNOR3X2_RVT




.subckt XOR2X1_RVT A1 A2 VDD VSS Y
MN7 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN5 Y1 A1B SA4 VSS n105 w=0.27u l=0.03u nf=1.0 m=1
MN4 SA2 A2B VSS VSS n105 w=0.23u l=0.03u nf=1.0 m=1
MN3 Y1 A1 SA2 VSS n105 w=0.23u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.21u l=0.03u nf=1.0 m=1
MN1 A1B A1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MP7 Y Y1 VDD VDD p105 w=0.75u l=0.03u nf=1.0 m=1
MP6 Y1 A1B SA3 VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.40u l=0.03u nf=1.0 m=1
MP4 Y1 A1 SA1 VDD p105 w=0.33u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.33u l=0.03u nf=1.0 m=1
MP2 A2B A2 VDD VDD p105 w=0.33u l=0.03u nf=1.0 m=1
MP1 A1B A1 VDD VDD p105 w=0.36u l=0.03u nf=1.0 m=1
.ends XOR2X1_RVT




.subckt XOR2X2_RVT A1 A2 VDD VSS Y
MP1 A1B A1 VDD VDD p105 w=0.63u l=0.03u nf=1.0 m=1
MP7 Y Y1 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP5 SA3 A2B VDD VDD p105 w=0.64u l=0.03u nf=1.0 m=1
MP4 Y1 A1 SA1 VDD p105 w=0.63u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.63u l=0.03u nf=1.0 m=1
MP2 A2B A2 VDD VDD p105 w=0.63u l=0.03u nf=1.0 m=1
MP6 Y1 A1B SA3 VDD p105 w=0.64u l=0.03u nf=1.0 m=1
MN4 SA2 A2B VSS VSS n105 w=0.40u l=0.03u nf=1.0 m=1
MN3 Y1 A1 SA2 VSS n105 w=0.40u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN1 A1B A1 VSS VSS n105 w=0.32u l=0.03u nf=1.0 m=1
MN7 Y Y1 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=2
MN6 SA4 A2 VSS VSS n105 w=0.38u l=0.03u nf=1.0 m=1
MN5 Y1 A1B SA4 VSS n105 w=0.38u l=0.03u nf=1.0 m=1
.ends XOR2X2_RVT




.subckt XOR3X1_RVT A1 A2 A3 VDD VSS Y
MP11 Y Y2 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=1
MP8 Y1B Y1 VDD VDD p105 w=0.37u l=0.03u nf=1.0 m=1
MP10 Y1 A3B Y2 VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP9 Y1B A3 Y2 VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.60u l=0.03u nf=1.0 m=2
MP7 A3B A3 VDD VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.55u l=0.03u nf=1.0 m=2
MP6 Y1 A1 SA3 VDD p105 w=0.60u l=0.03u nf=1.0 m=2
MP2 A2B A2 VDD VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MP4 Y1 A1B SA1 VDD p105 w=0.55u l=0.03u nf=1.0 m=2
MP1 A1B A1 VDD VDD p105 w=0.53u l=0.03u nf=1.0 m=1
MN11 Y Y2 VSS VSS n105 w=0.42u l=0.03u nf=1.0 m=1
MN8 Y1B Y1 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN10 Y1 A3 Y2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN9 Y1B A3B Y2 VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN1 A1B A1 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN5 Y1 A1 SA4 VSS n105 w=0.29u l=0.03u nf=1.0 m=2
MN4 SA2 A2B VSS VSS n105 w=0.25u l=0.03u nf=1.0 m=2
MN3 Y1 A1B SA2 VSS n105 w=0.25u l=0.03u nf=1.0 m=2
MN7 A3B A3 VSS VSS n105 w=0.3u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.29u l=0.03u nf=1.0 m=2
.ends XOR3X1_RVT




.subckt XOR3X2_RVT A1 A2 A3 VDD VSS Y
MP11 Y Y2 VDD VDD p105 w=0.8u l=0.03u nf=1.0 m=2
MP8 Y1B YA1 VDD VDD p105 w=0.80u l=0.03u nf=1.0 m=1
MP10 YA1 A3B Y2 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP9 Y1B A3 Y2 VDD p105 w=0.30u l=0.03u nf=1.0 m=1
MP5 SA3 A2B VDD VDD p105 w=0.70u l=0.03u nf=1.0 m=2
MP7 A3B A3 VDD VDD p105 w=0.45u l=0.03u nf=1.0 m=1
MP3 SA1 A2 VDD VDD p105 w=0.65u l=0.03u nf=1.0 m=2
MP6 YA1 A1 SA3 VDD p105 w=0.70u l=0.03u nf=1.0 m=2
MP2 A2B A2 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MP4 YA1 A1B SA1 VDD p105 w=0.65u l=0.03u nf=1.0 m=2
MP1 A1B A1 VDD VDD p105 w=0.39u l=0.03u nf=1.0 m=1
MN11 Y Y2 VSS VSS n105 w=0.40u l=0.03u nf=1.0 m=2
MN8 Y1B YA1 VSS VSS n105 w=0.35u l=0.03u nf=1.0 m=1
MN10 YA1 A3 Y2 VSS n105 w=0.30u l=0.03u nf=1.0 m=1
MN9 Y1B A3B Y2 VSS n105 w=0.30u l=0.03u nf=1.0 m=1
MN1 A1B A1 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN2 A2B A2 VSS VSS n105 w=0.20u l=0.03u nf=1.0 m=1
MN5 YA1 A1 SA4 VSS n105 w=0.28u l=0.03u nf=1.0 m=2
MN4 SA2 A2B VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=2
MN3 YA1 A1B SA2 VSS n105 w=0.28u l=0.03u nf=1.0 m=2
MN7 A3B A3 VSS VSS n105 w=0.15u l=0.03u nf=1.0 m=1
MN6 SA4 A2 VSS VSS n105 w=0.28u l=0.03u nf=1.0 m=2
.ends XOR3X2_RVT


