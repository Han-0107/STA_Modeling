* NAND Gate
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/SAED90nm/saed90nm.cdl
.include /data/yaohuihan/Research/STA_Modeling/gates/Libs/SAED90nm/SAED90nm.lib

.temp 25
.param VOL=1.1
VDD VDD 0 VOL
VSS VSS 0 0

VIN_AN an 0 PULSE(0 VOL 0 1.8n 1.8n 5n 40n)
VIN_B b 0 DC VOL

Cout y 0 0.1p

X1 an b y VDD VSS NAND2X1

.tran 0.000001n 10n

.measure tran tpHL TRIG V(an) VAL=0.55 FALL=1 TARG V(y) VAL=0.55 RISE=1
.measure tran tpLH TRIG V(an) VAL=0.55 RISE=1 TARG V(y) VAL=0.55 FALL=1

.end
